VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO collatz
  CLASS BLOCK ;
  FOREIGN collatz ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.000 BY 220.000 ;
  PIN bs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 216.000 109.760 220.000 110.320 ;
    END
  END bs
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END clk
  PIN co[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 5.600 0.000 6.160 4.000 ;
    END
  END co[0]
  PIN co[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END co[10]
  PIN co[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END co[11]
  PIN co[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END co[12]
  PIN co[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END co[13]
  PIN co[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END co[14]
  PIN co[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END co[15]
  PIN co[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 0.000 12.880 4.000 ;
    END
  END co[1]
  PIN co[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 4.000 ;
    END
  END co[2]
  PIN co[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END co[3]
  PIN co[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END co[4]
  PIN co[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 4.000 ;
    END
  END co[5]
  PIN co[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END co[6]
  PIN co[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END co[7]
  PIN co[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END co[8]
  PIN co[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END co[9]
  PIN st
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END st
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 204.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 204.140 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 204.140 ;
    END
  END vss
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 4.000 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END x[11]
  PIN x[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END x[12]
  PIN x[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END x[13]
  PIN x[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END x[14]
  PIN x[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END x[15]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END x[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 212.800 204.140 ;
      LAYER Metal2 ;
        RECT 5.180 4.300 214.900 204.030 ;
        RECT 5.180 3.500 5.300 4.300 ;
        RECT 6.460 3.500 12.020 4.300 ;
        RECT 13.180 3.500 18.740 4.300 ;
        RECT 19.900 3.500 25.460 4.300 ;
        RECT 26.620 3.500 32.180 4.300 ;
        RECT 33.340 3.500 38.900 4.300 ;
        RECT 40.060 3.500 45.620 4.300 ;
        RECT 46.780 3.500 52.340 4.300 ;
        RECT 53.500 3.500 59.060 4.300 ;
        RECT 60.220 3.500 65.780 4.300 ;
        RECT 66.940 3.500 72.500 4.300 ;
        RECT 73.660 3.500 79.220 4.300 ;
        RECT 80.380 3.500 85.940 4.300 ;
        RECT 87.100 3.500 92.660 4.300 ;
        RECT 93.820 3.500 99.380 4.300 ;
        RECT 100.540 3.500 106.100 4.300 ;
        RECT 107.260 3.500 112.820 4.300 ;
        RECT 113.980 3.500 119.540 4.300 ;
        RECT 120.700 3.500 126.260 4.300 ;
        RECT 127.420 3.500 132.980 4.300 ;
        RECT 134.140 3.500 139.700 4.300 ;
        RECT 140.860 3.500 146.420 4.300 ;
        RECT 147.580 3.500 153.140 4.300 ;
        RECT 154.300 3.500 159.860 4.300 ;
        RECT 161.020 3.500 166.580 4.300 ;
        RECT 167.740 3.500 173.300 4.300 ;
        RECT 174.460 3.500 180.020 4.300 ;
        RECT 181.180 3.500 186.740 4.300 ;
        RECT 187.900 3.500 193.460 4.300 ;
        RECT 194.620 3.500 200.180 4.300 ;
        RECT 201.340 3.500 206.900 4.300 ;
        RECT 208.060 3.500 213.620 4.300 ;
        RECT 214.780 3.500 214.900 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 165.500 216.000 203.980 ;
        RECT 4.300 164.340 216.000 165.500 ;
        RECT 3.500 110.620 216.000 164.340 ;
        RECT 3.500 109.460 215.700 110.620 ;
        RECT 3.500 55.740 216.000 109.460 ;
        RECT 4.300 54.580 216.000 55.740 ;
        RECT 3.500 12.460 216.000 54.580 ;
      LAYER Metal4 ;
        RECT 9.100 15.080 21.940 127.590 ;
        RECT 24.140 15.080 98.740 127.590 ;
        RECT 100.940 15.080 175.540 127.590 ;
        RECT 177.740 15.080 193.060 127.590 ;
        RECT 9.100 14.650 193.060 15.080 ;
  END
END collatz
END LIBRARY

