// This is the unpowered netlist.
module collatz (bs,
    clk,
    st,
    co,
    x);
 output bs;
 input clk;
 input st;
 input [15:0] co;
 output [15:0] x;

 wire \Datapath.i[0] ;
 wire \Datapath.i[10] ;
 wire \Datapath.i[11] ;
 wire \Datapath.i[12] ;
 wire \Datapath.i[13] ;
 wire \Datapath.i[14] ;
 wire \Datapath.i[15] ;
 wire \Datapath.i[1] ;
 wire \Datapath.i[2] ;
 wire \Datapath.i[3] ;
 wire \Datapath.i[4] ;
 wire \Datapath.i[5] ;
 wire \Datapath.i[6] ;
 wire \Datapath.i[7] ;
 wire \Datapath.i[8] ;
 wire \Datapath.i[9] ;
 wire \Datapath.k[0] ;
 wire \Datapath.k[10] ;
 wire \Datapath.k[11] ;
 wire \Datapath.k[12] ;
 wire \Datapath.k[13] ;
 wire \Datapath.k[14] ;
 wire \Datapath.k[15] ;
 wire \Datapath.k[16] ;
 wire \Datapath.k[17] ;
 wire \Datapath.k[18] ;
 wire \Datapath.k[19] ;
 wire \Datapath.k[1] ;
 wire \Datapath.k[2] ;
 wire \Datapath.k[3] ;
 wire \Datapath.k[4] ;
 wire \Datapath.k[5] ;
 wire \Datapath.k[6] ;
 wire \Datapath.k[7] ;
 wire \Datapath.k[8] ;
 wire \Datapath.k[9] ;
 wire \FSM.CS[0] ;
 wire \FSM.CS[1] ;
 wire \FSM.NS[0] ;
 wire \FSM.NS[1] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _344_ (.I(\FSM.CS[0] ),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _345_ (.I(\FSM.CS[1] ),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _346_ (.I(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _347_ (.A1(_036_),
    .A2(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _348_ (.I(_039_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _349_ (.I(\Datapath.i[0] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _350_ (.A1(net18),
    .A2(_040_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _351_ (.I(_039_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _352_ (.I(_041_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _353_ (.A1(_042_),
    .A2(\Datapath.i[1] ),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _354_ (.I(_043_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _355_ (.A1(_042_),
    .A2(\Datapath.i[2] ),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _356_ (.I(_044_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _357_ (.I(\Datapath.i[3] ),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _358_ (.A1(net18),
    .A2(_045_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _359_ (.I(_041_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _360_ (.I(_046_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _361_ (.A1(_047_),
    .A2(\Datapath.i[4] ),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _362_ (.I(_048_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _363_ (.A1(_047_),
    .A2(\Datapath.i[5] ),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _364_ (.I(_049_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _365_ (.I(\Datapath.i[6] ),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _366_ (.A1(net18),
    .A2(_050_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _367_ (.I(\Datapath.i[7] ),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _368_ (.A1(net18),
    .A2(_051_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _369_ (.I(\Datapath.i[8] ),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _370_ (.A1(net18),
    .A2(_052_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _371_ (.I(\Datapath.i[9] ),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _372_ (.A1(net18),
    .A2(_053_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _373_ (.A1(_047_),
    .A2(\Datapath.i[10] ),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _374_ (.I(_054_),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _375_ (.I(\Datapath.i[11] ),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _376_ (.A1(net18),
    .A2(_055_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _377_ (.I(\Datapath.i[12] ),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _378_ (.A1(net18),
    .A2(_056_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _379_ (.I(\Datapath.i[13] ),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _380_ (.A1(net18),
    .A2(_057_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _381_ (.I(\Datapath.i[14] ),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _382_ (.A1(_039_),
    .A2(_058_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _383_ (.I(\Datapath.i[15] ),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _384_ (.A1(_039_),
    .A2(_059_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _385_ (.I(\FSM.CS[0] ),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _386_ (.A1(_038_),
    .A2(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _387_ (.I(_061_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _388_ (.A1(_047_),
    .A2(net17),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _389_ (.I(_036_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _390_ (.I(\Datapath.k[1] ),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _391_ (.A1(_064_),
    .A2(_065_),
    .B(_037_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _392_ (.A1(net1),
    .A2(_062_),
    .B(_063_),
    .C(_066_),
    .ZN(\FSM.NS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _393_ (.A1(net16),
    .A2(net2),
    .A3(net3),
    .A4(net4),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _394_ (.A1(net12),
    .A2(net13),
    .A3(net14),
    .A4(net15),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _395_ (.A1(_067_),
    .A2(_068_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _396_ (.A1(_069_),
    .A2(net5),
    .A3(net6),
    .A4(net7),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _397_ (.A1(net8),
    .A2(net9),
    .A3(net10),
    .A4(net11),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _398_ (.A1(_070_),
    .A2(_060_),
    .A3(net1),
    .A4(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _399_ (.A1(_060_),
    .A2(_037_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _400_ (.A1(_072_),
    .A2(_039_),
    .A3(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _401_ (.I(\Datapath.k[9] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _402_ (.I(\Datapath.k[8] ),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _403_ (.A1(_075_),
    .A2(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _404_ (.A1(\Datapath.k[19] ),
    .A2(\Datapath.k[18] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _405_ (.I(\Datapath.k[11] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _406_ (.I(\Datapath.k[10] ),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _407_ (.A1(_079_),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _408_ (.I(\Datapath.k[17] ),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _409_ (.I(\Datapath.k[16] ),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _410_ (.A1(_082_),
    .A2(_083_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _411_ (.A1(_077_),
    .A2(_078_),
    .A3(_081_),
    .A4(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _412_ (.I(\Datapath.k[0] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _413_ (.A1(\Datapath.k[5] ),
    .A2(\Datapath.k[4] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _414_ (.I(\Datapath.k[15] ),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _415_ (.I(\Datapath.k[14] ),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _416_ (.A1(_088_),
    .A2(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _417_ (.I(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _418_ (.A1(_085_),
    .A2(_086_),
    .A3(_087_),
    .A4(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _419_ (.A1(\Datapath.k[7] ),
    .A2(\Datapath.k[6] ),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _420_ (.I(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _421_ (.I(\Datapath.k[3] ),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _422_ (.I(\Datapath.k[2] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _423_ (.A1(_095_),
    .A2(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _424_ (.I(\Datapath.k[13] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _425_ (.I(\Datapath.k[12] ),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _426_ (.A1(_098_),
    .A2(_099_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _427_ (.A1(_065_),
    .A2(_094_),
    .A3(_097_),
    .A4(_100_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _428_ (.I(_073_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _429_ (.I(_102_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _430_ (.A1(_092_),
    .A2(_101_),
    .B(_103_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _431_ (.A1(_074_),
    .A2(_104_),
    .ZN(\FSM.NS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _432_ (.A1(_040_),
    .A2(_037_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _433_ (.A1(_039_),
    .A2(_040_),
    .B(_105_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _434_ (.A1(\Datapath.i[1] ),
    .A2(\Datapath.i[0] ),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _435_ (.A1(_106_),
    .A2(_037_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _436_ (.I(\Datapath.i[1] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _437_ (.A1(_043_),
    .A2(_107_),
    .B1(_108_),
    .B2(_040_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _438_ (.I(\Datapath.i[2] ),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _439_ (.A1(_106_),
    .A2(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _440_ (.I(_110_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _441_ (.A1(_111_),
    .A2(_037_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _442_ (.A1(_112_),
    .A2(_044_),
    .B1(_109_),
    .B2(_106_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _443_ (.A1(_110_),
    .A2(_037_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _444_ (.A1(_062_),
    .A2(\Datapath.i[3] ),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _445_ (.A1(_113_),
    .A2(_045_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _446_ (.A1(_113_),
    .A2(_114_),
    .B(_115_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _447_ (.A1(_115_),
    .A2(\Datapath.i[4] ),
    .B(_062_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _448_ (.A1(_115_),
    .A2(\Datapath.i[4] ),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _449_ (.I(_117_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _450_ (.A1(_116_),
    .A2(_118_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _451_ (.A1(_118_),
    .A2(\Datapath.i[5] ),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _452_ (.I(_061_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _453_ (.I(_120_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _454_ (.A1(\Datapath.i[5] ),
    .A2(\Datapath.i[4] ),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _455_ (.A1(_122_),
    .A2(_045_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _456_ (.I(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _457_ (.A1(_113_),
    .A2(_124_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _458_ (.A1(_119_),
    .A2(_121_),
    .A3(_125_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _459_ (.A1(_125_),
    .A2(\Datapath.i[6] ),
    .B(_062_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _460_ (.A1(_125_),
    .A2(\Datapath.i[6] ),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _461_ (.I(_127_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _462_ (.A1(_126_),
    .A2(_128_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _463_ (.A1(_128_),
    .A2(\Datapath.i[7] ),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _464_ (.A1(_129_),
    .A2(_062_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _465_ (.A1(_051_),
    .A2(_127_),
    .B(_130_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _466_ (.A1(_128_),
    .A2(\Datapath.i[8] ),
    .A3(\Datapath.i[7] ),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _467_ (.A1(_131_),
    .A2(_062_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _468_ (.A1(_052_),
    .A2(_129_),
    .B(_132_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _469_ (.A1(_131_),
    .A2(_053_),
    .B(_062_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _470_ (.A1(_053_),
    .A2(_131_),
    .B(_133_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _471_ (.A1(_062_),
    .A2(\Datapath.i[10] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _472_ (.A1(_111_),
    .A2(_051_),
    .A3(_050_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _473_ (.A1(\Datapath.i[9] ),
    .A2(\Datapath.i[8] ),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _474_ (.I(_136_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _475_ (.A1(_135_),
    .A2(_037_),
    .A3(_123_),
    .A4(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _476_ (.I(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _477_ (.A1(_139_),
    .A2(\Datapath.i[10] ),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _478_ (.I(_140_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _479_ (.A1(_134_),
    .A2(_138_),
    .B(_141_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _480_ (.A1(_131_),
    .A2(_053_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _481_ (.A1(_142_),
    .A2(\Datapath.i[11] ),
    .A3(\Datapath.i[10] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _482_ (.A1(_143_),
    .A2(_062_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _483_ (.A1(_055_),
    .A2(_140_),
    .B(_144_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _484_ (.A1(_141_),
    .A2(\Datapath.i[11] ),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _485_ (.A1(_143_),
    .A2(_056_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _486_ (.I(_146_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _487_ (.A1(_147_),
    .A2(_062_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _488_ (.A1(_056_),
    .A2(_145_),
    .B(_148_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _489_ (.A1(_141_),
    .A2(\Datapath.i[13] ),
    .A3(\Datapath.i[12] ),
    .A4(\Datapath.i[11] ),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _490_ (.A1(\Datapath.i[13] ),
    .A2(_146_),
    .B(_149_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _491_ (.A1(_150_),
    .A2(_121_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _492_ (.A1(_149_),
    .A2(_058_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _493_ (.A1(_149_),
    .A2(_058_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _494_ (.A1(_151_),
    .A2(_152_),
    .A3(_121_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _495_ (.A1(_152_),
    .A2(\Datapath.i[15] ),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _496_ (.A1(_149_),
    .A2(_059_),
    .A3(_058_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _497_ (.A1(_153_),
    .A2(_154_),
    .A3(_121_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _498_ (.A1(_060_),
    .A2(\Datapath.k[0] ),
    .B(_037_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _499_ (.A1(_064_),
    .A2(net1),
    .B(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _500_ (.A1(_103_),
    .A2(\Datapath.k[1] ),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _501_ (.I(_042_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _502_ (.A1(_156_),
    .A2(_157_),
    .B1(_086_),
    .B2(_158_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _503_ (.A1(_121_),
    .A2(net8),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _504_ (.A1(_060_),
    .A2(_065_),
    .B1(_096_),
    .B2(_073_),
    .C(_159_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _505_ (.A1(net9),
    .A2(_121_),
    .B1(\Datapath.k[3] ),
    .B2(_103_),
    .C(_042_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _506_ (.A1(_096_),
    .A2(_065_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _507_ (.A1(\Datapath.k[2] ),
    .A2(\Datapath.k[1] ),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _508_ (.A1(_161_),
    .A2(_162_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _509_ (.A1(_163_),
    .A2(_086_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _510_ (.A1(_161_),
    .A2(\Datapath.k[0] ),
    .A3(_162_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _511_ (.A1(_164_),
    .A2(_036_),
    .A3(_165_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _512_ (.A1(_160_),
    .A2(_166_),
    .B1(_096_),
    .B2(_158_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _513_ (.A1(_165_),
    .A2(_162_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _514_ (.A1(\Datapath.k[3] ),
    .A2(\Datapath.k[2] ),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _515_ (.A1(_167_),
    .A2(_097_),
    .A3(_168_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _516_ (.A1(_097_),
    .A2(_168_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _517_ (.A1(_165_),
    .A2(_162_),
    .A3(_170_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _518_ (.A1(_169_),
    .A2(_064_),
    .A3(_171_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _519_ (.A1(net10),
    .A2(_121_),
    .B1(\Datapath.k[4] ),
    .B2(_102_),
    .C(_042_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _520_ (.A1(_172_),
    .A2(_173_),
    .B1(_095_),
    .B2(_158_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _521_ (.A1(\Datapath.k[3] ),
    .A2(\Datapath.k[1] ),
    .B(\Datapath.k[2] ),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _522_ (.A1(_165_),
    .A2(_170_),
    .B(_174_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _523_ (.A1(\Datapath.k[4] ),
    .A2(\Datapath.k[3] ),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _524_ (.I(_176_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _525_ (.A1(\Datapath.k[4] ),
    .A2(\Datapath.k[3] ),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _526_ (.A1(_177_),
    .A2(_178_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _527_ (.A1(_175_),
    .A2(_179_),
    .Z(_180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _528_ (.A1(_175_),
    .A2(_179_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _529_ (.A1(_180_),
    .A2(_064_),
    .A3(_181_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _530_ (.A1(net11),
    .A2(_120_),
    .B1(\Datapath.k[5] ),
    .B2(_102_),
    .C(_042_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _531_ (.I(\Datapath.k[4] ),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _532_ (.A1(_182_),
    .A2(_183_),
    .B1(_184_),
    .B2(_158_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _533_ (.A1(_181_),
    .A2(_176_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _534_ (.I(\Datapath.k[5] ),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _535_ (.A1(_186_),
    .A2(_184_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _536_ (.A1(_187_),
    .A2(_087_),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _537_ (.A1(_185_),
    .A2(_188_),
    .B(_060_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _538_ (.A1(_185_),
    .A2(_188_),
    .B(_189_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _539_ (.A1(net12),
    .A2(_120_),
    .B1(\Datapath.k[6] ),
    .B2(_102_),
    .C(_042_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _540_ (.A1(_190_),
    .A2(_191_),
    .B1(_186_),
    .B2(_158_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _541_ (.A1(_186_),
    .A2(_095_),
    .B(_184_),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _542_ (.I(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _543_ (.A1(_181_),
    .A2(_193_),
    .B(_087_),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _544_ (.A1(\Datapath.k[6] ),
    .A2(\Datapath.k[5] ),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _545_ (.I(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _546_ (.A1(\Datapath.k[6] ),
    .A2(\Datapath.k[5] ),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _547_ (.A1(_196_),
    .A2(_197_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _548_ (.A1(_194_),
    .A2(_198_),
    .Z(_199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _549_ (.A1(_194_),
    .A2(_198_),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _550_ (.A1(_199_),
    .A2(_200_),
    .A3(_036_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _551_ (.A1(net13),
    .A2(_120_),
    .B1(\Datapath.k[7] ),
    .B2(_102_),
    .C(_046_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _552_ (.I(\Datapath.k[6] ),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _553_ (.A1(_201_),
    .A2(_202_),
    .B1(_203_),
    .B2(_158_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _554_ (.A1(_200_),
    .A2(_195_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _555_ (.A1(\Datapath.k[7] ),
    .A2(\Datapath.k[6] ),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _556_ (.I(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _557_ (.A1(_206_),
    .A2(_093_),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _558_ (.A1(_204_),
    .A2(_207_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _559_ (.A1(_094_),
    .A2(_205_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _560_ (.A1(_200_),
    .A2(_195_),
    .A3(_209_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _561_ (.A1(_208_),
    .A2(_064_),
    .A3(_210_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _562_ (.A1(net14),
    .A2(_120_),
    .B1(\Datapath.k[8] ),
    .B2(_102_),
    .C(_046_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _563_ (.I(\Datapath.k[7] ),
    .ZN(_213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _564_ (.A1(_211_),
    .A2(_212_),
    .B1(_213_),
    .B2(_158_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _565_ (.A1(_188_),
    .A2(_179_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _566_ (.A1(_198_),
    .A2(_207_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _567_ (.A1(_214_),
    .A2(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _568_ (.A1(_175_),
    .A2(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _569_ (.I(_215_),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _570_ (.A1(_195_),
    .A2(_205_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _571_ (.A1(_218_),
    .A2(_192_),
    .B(_219_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _572_ (.A1(_217_),
    .A2(_220_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _573_ (.I(_221_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _574_ (.A1(_076_),
    .A2(_213_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _575_ (.A1(\Datapath.k[8] ),
    .A2(\Datapath.k[7] ),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _576_ (.A1(_223_),
    .A2(_224_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _577_ (.A1(_222_),
    .A2(_225_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _578_ (.I(_226_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _579_ (.A1(_222_),
    .A2(_225_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _580_ (.A1(_227_),
    .A2(_064_),
    .A3(_228_),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _581_ (.A1(net15),
    .A2(_120_),
    .B1(\Datapath.k[9] ),
    .B2(_102_),
    .C(_046_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _582_ (.A1(_229_),
    .A2(_230_),
    .B1(_076_),
    .B2(_158_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _583_ (.A1(_227_),
    .A2(_224_),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _584_ (.A1(\Datapath.k[9] ),
    .A2(\Datapath.k[8] ),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _585_ (.A1(_077_),
    .A2(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _586_ (.I(_233_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _587_ (.A1(_231_),
    .A2(_234_),
    .B(_060_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _588_ (.A1(_231_),
    .A2(_234_),
    .B(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _589_ (.A1(\Datapath.k[10] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net16),
    .C(_046_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _590_ (.A1(_236_),
    .A2(_237_),
    .B1(_075_),
    .B2(_158_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _591_ (.A1(_225_),
    .A2(_233_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _592_ (.A1(_224_),
    .A2(_232_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _593_ (.A1(_221_),
    .A2(_238_),
    .B(_239_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _594_ (.A1(_080_),
    .A2(_075_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _595_ (.A1(\Datapath.k[10] ),
    .A2(\Datapath.k[9] ),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _596_ (.A1(_241_),
    .A2(_242_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _597_ (.A1(_240_),
    .A2(_243_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _598_ (.A1(_240_),
    .A2(_243_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _599_ (.A1(_244_),
    .A2(_064_),
    .A3(_245_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _600_ (.A1(\Datapath.k[11] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net2),
    .C(_046_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _601_ (.A1(_246_),
    .A2(_247_),
    .B1(_080_),
    .B2(_158_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _602_ (.A1(\Datapath.k[11] ),
    .A2(\Datapath.k[10] ),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _603_ (.A1(_081_),
    .A2(_248_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _604_ (.A1(_244_),
    .A2(_242_),
    .A3(_249_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _605_ (.A1(_250_),
    .A2(_036_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _606_ (.A1(_244_),
    .A2(_242_),
    .B(_249_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _607_ (.A1(_251_),
    .A2(_252_),
    .Z(_253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _608_ (.A1(\Datapath.k[12] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net3),
    .C(_046_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _609_ (.A1(_253_),
    .A2(_254_),
    .B1(_079_),
    .B2(_047_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _610_ (.A1(_243_),
    .A2(_249_),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _611_ (.A1(_238_),
    .A2(_255_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _612_ (.A1(_217_),
    .A2(_220_),
    .B(_256_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _613_ (.A1(_255_),
    .A2(_239_),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _614_ (.A1(_258_),
    .A2(_242_),
    .A3(_248_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _615_ (.A1(_257_),
    .A2(_259_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _616_ (.I(_260_),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _617_ (.A1(_099_),
    .A2(_079_),
    .ZN(_262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _618_ (.A1(\Datapath.k[12] ),
    .A2(\Datapath.k[11] ),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _619_ (.A1(_261_),
    .A2(_262_),
    .A3(_263_),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _620_ (.A1(_262_),
    .A2(_263_),
    .ZN(_265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _621_ (.A1(_260_),
    .A2(_265_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _622_ (.A1(_264_),
    .A2(_064_),
    .A3(_266_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _623_ (.A1(\Datapath.k[13] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net4),
    .C(_046_),
    .ZN(_268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _624_ (.A1(_267_),
    .A2(_268_),
    .B1(_099_),
    .B2(_047_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _625_ (.I(_263_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _626_ (.A1(_261_),
    .A2(_262_),
    .B(_269_),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _627_ (.A1(\Datapath.k[13] ),
    .A2(\Datapath.k[12] ),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _628_ (.A1(_100_),
    .A2(_271_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _629_ (.A1(_270_),
    .A2(_272_),
    .Z(_273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _630_ (.A1(_270_),
    .A2(_272_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _631_ (.A1(_273_),
    .A2(_274_),
    .A3(_036_),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _632_ (.A1(\Datapath.k[14] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net5),
    .C(_046_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _633_ (.A1(_275_),
    .A2(_276_),
    .B1(_098_),
    .B2(_047_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _634_ (.A1(_265_),
    .A2(_272_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _635_ (.A1(_257_),
    .A2(_259_),
    .B(_277_),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _636_ (.A1(_263_),
    .A2(_271_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _637_ (.I(_279_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _638_ (.A1(_278_),
    .A2(_280_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _639_ (.A1(_089_),
    .A2(_098_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _640_ (.A1(\Datapath.k[14] ),
    .A2(\Datapath.k[13] ),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _641_ (.A1(_282_),
    .A2(_283_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _642_ (.I(_284_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _643_ (.A1(_281_),
    .A2(_285_),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _644_ (.A1(_278_),
    .A2(_280_),
    .A3(_284_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _645_ (.A1(_286_),
    .A2(_064_),
    .A3(_287_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _646_ (.A1(\Datapath.k[15] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net6),
    .C(_046_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _647_ (.A1(_288_),
    .A2(_289_),
    .B1(_089_),
    .B2(_047_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _648_ (.A1(_278_),
    .A2(_280_),
    .B(_284_),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _649_ (.I(_283_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _650_ (.A1(\Datapath.k[15] ),
    .A2(\Datapath.k[14] ),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _651_ (.A1(_090_),
    .A2(_292_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _652_ (.I(_293_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _653_ (.A1(_290_),
    .A2(_291_),
    .B(_294_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _654_ (.A1(_286_),
    .A2(_283_),
    .A3(_293_),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _655_ (.A1(_295_),
    .A2(_296_),
    .A3(_064_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _656_ (.A1(\Datapath.k[16] ),
    .A2(_103_),
    .B1(_038_),
    .B2(net7),
    .C(_042_),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _657_ (.A1(_039_),
    .A2(\Datapath.k[15] ),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _658_ (.A1(_297_),
    .A2(_298_),
    .B(_299_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _659_ (.A1(_284_),
    .A2(_293_),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _660_ (.A1(_277_),
    .A2(_300_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _661_ (.I(_301_),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _662_ (.A1(_302_),
    .A2(_238_),
    .A3(_255_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _663_ (.A1(_222_),
    .A2(_303_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _664_ (.A1(_259_),
    .A2(_302_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _665_ (.A1(_283_),
    .A2(_292_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _666_ (.A1(_300_),
    .A2(_279_),
    .B(_306_),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _667_ (.A1(_305_),
    .A2(_307_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _668_ (.A1(_304_),
    .A2(_308_),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _669_ (.A1(_083_),
    .A2(_088_),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _670_ (.A1(\Datapath.k[16] ),
    .A2(\Datapath.k[15] ),
    .ZN(_311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _671_ (.A1(_310_),
    .A2(_311_),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _672_ (.A1(_309_),
    .A2(_312_),
    .ZN(_313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _673_ (.I(_312_),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _674_ (.A1(_304_),
    .A2(_308_),
    .B(_314_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _675_ (.A1(_036_),
    .A2(_037_),
    .ZN(_316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _676_ (.I(_316_),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _677_ (.A1(_313_),
    .A2(_315_),
    .A3(_317_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _678_ (.A1(_047_),
    .A2(\Datapath.k[16] ),
    .B1(\Datapath.k[17] ),
    .B2(_060_),
    .ZN(_319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _679_ (.A1(_318_),
    .A2(_319_),
    .B(_121_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _680_ (.A1(_315_),
    .A2(_311_),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _681_ (.A1(\Datapath.k[17] ),
    .A2(\Datapath.k[16] ),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _682_ (.A1(_320_),
    .A2(_084_),
    .A3(_321_),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _683_ (.A1(_084_),
    .A2(_321_),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _684_ (.A1(_315_),
    .A2(_311_),
    .A3(_323_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _685_ (.A1(_322_),
    .A2(_317_),
    .A3(_324_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _686_ (.A1(_042_),
    .A2(\Datapath.k[17] ),
    .B1(\Datapath.k[18] ),
    .B2(_060_),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _687_ (.A1(_325_),
    .A2(_326_),
    .B(_121_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _688_ (.A1(_314_),
    .A2(_084_),
    .A3(_321_),
    .ZN(_327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _689_ (.A1(\Datapath.k[17] ),
    .A2(\Datapath.k[15] ),
    .B(\Datapath.k[16] ),
    .ZN(_328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _690_ (.A1(_309_),
    .A2(_327_),
    .B(_328_),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _691_ (.A1(\Datapath.k[18] ),
    .A2(\Datapath.k[17] ),
    .Z(_330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _692_ (.A1(\Datapath.k[18] ),
    .A2(\Datapath.k[17] ),
    .ZN(_331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _693_ (.A1(_330_),
    .A2(_331_),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _694_ (.I(_332_),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _695_ (.A1(_329_),
    .A2(_333_),
    .Z(_334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _696_ (.A1(_329_),
    .A2(_333_),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _697_ (.A1(_334_),
    .A2(_317_),
    .A3(_335_),
    .ZN(_336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _698_ (.A1(_042_),
    .A2(\Datapath.k[18] ),
    .B1(\Datapath.k[19] ),
    .B2(_060_),
    .ZN(_337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _699_ (.A1(_336_),
    .A2(_337_),
    .B(_121_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _700_ (.A1(\Datapath.k[19] ),
    .A2(\Datapath.k[18] ),
    .ZN(_338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _701_ (.A1(_078_),
    .A2(_338_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _702_ (.A1(_335_),
    .A2(_331_),
    .A3(_339_),
    .ZN(_340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _703_ (.A1(_340_),
    .A2(_317_),
    .ZN(_341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _704_ (.A1(_335_),
    .A2(_331_),
    .B(_339_),
    .ZN(_342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _705_ (.A1(_047_),
    .A2(\Datapath.k[19] ),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _706_ (.A1(_341_),
    .A2(_342_),
    .B(_343_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _707_ (.D(_000_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _708_ (.D(_001_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _709_ (.D(_002_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _710_ (.D(_003_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _711_ (.D(_004_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _712_ (.D(_005_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _713_ (.D(_006_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _714_ (.D(_007_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _715_ (.D(_008_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _716_ (.D(_009_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _717_ (.D(_010_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _718_ (.D(_011_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _719_ (.D(_012_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _720_ (.D(_013_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _721_ (.D(_014_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _722_ (.D(_015_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _723_ (.D(_016_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _724_ (.D(_017_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _725_ (.D(_018_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _726_ (.D(_019_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _727_ (.D(_020_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _728_ (.D(_021_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _729_ (.D(_022_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _730_ (.D(_023_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _731_ (.D(_024_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _732_ (.D(_025_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _733_ (.D(_026_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _734_ (.D(_027_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _735_ (.D(_028_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _736_ (.D(_029_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _737_ (.D(_030_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _738_ (.D(_031_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _739_ (.D(_032_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _740_ (.D(_033_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _741_ (.D(_034_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _742_ (.D(_035_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _743_ (.D(\FSM.NS[0] ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\FSM.CS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _744_ (.D(\FSM.NS[1] ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input1 (.I(co[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(co[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(co[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(co[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(co[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(co[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(co[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(co[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(co[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(co[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(co[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(co[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(co[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(co[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(co[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(co[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(st),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(bs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(x[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(x[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(x[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(x[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(x[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(x[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(x[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(x[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(x[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(x[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(x[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(x[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(x[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(x[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(x[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(x[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__A2 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__I (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A3 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__A2 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__A2 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A2 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A4 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__A2 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A2 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__I (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A2 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A2 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A2 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A2 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A1 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A2 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__A2 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A3 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A2 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__I (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A2 (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A2 (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__I (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A1 (.I(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__I (.I(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__618__A2 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__602__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__I (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__627__A2 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__618__A1 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__A1 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__I (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__A2 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__670__A2 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__A2 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__650__A1 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__A1 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__I (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__B (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__681__A2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__A2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__670__A1 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__A1 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__I (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__692__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__691__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__681__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__B1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__I (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__I (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__B (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__A2 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__A1 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__I (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__A2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__B1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__I (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__I (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__A1 (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A1 (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__B1 (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A2 (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A2 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__A2 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__I (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__B1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__552__I (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__A1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__B1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__A2 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__I (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__B1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__A2 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__A1 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__B1 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__I (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__595__A2 (.I(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__A1 (.I(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__B1 (.I(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__I (.I(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__631__A3 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__605__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__A3 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__I (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__B (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__B (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__I (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__B1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A2 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__I (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__B2 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A2 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__A2 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__698__A1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__A1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__C (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__C (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__C (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__C (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__C (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__I (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__A1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__A1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__C (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__I (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__705__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__B2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__633__B2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__624__B2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__609__B2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A1 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__A2 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A1 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__A2 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A2 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__A2 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__A2 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__488__A1 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__698__B2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__B2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__B2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__B (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__B (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__I (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__I (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__B (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__467__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__B (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__B (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__655__A3 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__645__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__622__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__599__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__A1 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A2 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__B1 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A1 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__B1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__701__A1 (.I(_078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A2 (.I(_078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__617__A2 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__609__B1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__603__A1 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A3 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__651__A1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__417__I (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__A2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__I (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A1 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A2 (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__B1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__B1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A2 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__A1 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__A2 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A3 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__A1 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A4 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__B2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__I (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__608__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__A2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__B2 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__A1 (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__B (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__699__B (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__687__B (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__679__B (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A1 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A3 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A2 (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A1 (.I(_128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A1 (.I(_128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__A2 (.I(_128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A2 (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A1 (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A1 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__469__A1 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__467__A1 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__479__A2 (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__I (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A1 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__A1 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__479__B (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A1 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A1 (.I(_143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__A1 (.I(_143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__A2 (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__486__I (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__487__A1 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__601__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__B2 (.I(_158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__C (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A2 (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__A2 (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__A3 (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A2 (.I(_162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__A1 (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A1 (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__A1 (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A3 (.I(_165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__A2 (.I(_168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__A3 (.I(_168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__A2 (.I(_170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A3 (.I(_170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__A1 (.I(_175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A1 (.I(_175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__A1 (.I(_175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__A2 (.I(_176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__I (.I(_176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__A2 (.I(_178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__565__A2 (.I(_179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__A2 (.I(_179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__A2 (.I(_179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__A1 (.I(_181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__A1 (.I(_181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A3 (.I(_181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__B (.I(_184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__A2 (.I(_184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__B1 (.I(_184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__A1 (.I(_185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__A1 (.I(_185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__A1 (.I(_186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B1 (.I(_186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__A1 (.I(_186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__565__A1 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__A2 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__A2 (.I(_188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__549__A1 (.I(_194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__A1 (.I(_194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__A1 (.I(_195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A2 (.I(_195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__A2 (.I(_195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__I (.I(_195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__A1 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__549__A2 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__A2 (.I(_198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A1 (.I(_200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__A1 (.I(_200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__A2 (.I(_200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__B1 (.I(_203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__558__A1 (.I(_204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__A2 (.I(_205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A2 (.I(_205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__I (.I(_205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__A1 (.I(_206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__566__A2 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__558__A2 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A3 (.I(_209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__A2 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B1 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A1 (.I(_214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__I (.I(_215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A2 (.I(_215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__612__A1 (.I(_217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__A1 (.I(_217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__571__B (.I(_219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__612__A2 (.I(_220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__A2 (.I(_220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__I (.I(_226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A1 (.I(_231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__A1 (.I(_231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__591__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__586__I (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A2 (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__A2 (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__658__A1 (.I(_297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__674__A1 (.I(_304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__668__A1 (.I(_304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__674__A2 (.I(_308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__668__A2 (.I(_308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(co[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(co[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(co[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(co[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(co[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(co[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(co[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(co[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(co[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(co[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(co[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(co[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(co[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(co[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(co[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(co[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(st));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A3 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__623__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__A4 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__632__B2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__646__B2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A3 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__B2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A4 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__380__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__372__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__708__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__714__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__715__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__717__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__718__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__722__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__711__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__712__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__721__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__724__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__744__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__719__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__720__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__725__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__726__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__727__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__728__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__730__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__731__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__733__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__723__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__735__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__736__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__738__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__739__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__740__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__741__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__742__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
endmodule

