magic
tech gf180mcuC
magscale 1 10
timestamp 1670102149
<< metal1 >>
rect 7074 77646 7086 77698
rect 7138 77695 7150 77698
rect 9650 77695 9662 77698
rect 7138 77649 9662 77695
rect 7138 77646 7150 77649
rect 9650 77646 9662 77649
rect 9714 77646 9726 77698
rect 11778 76974 11790 77026
rect 11842 77023 11854 77026
rect 12338 77023 12350 77026
rect 11842 76977 12350 77023
rect 11842 76974 11854 76977
rect 12338 76974 12350 76977
rect 12402 76974 12414 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 2046 76690 2098 76702
rect 2046 76626 2098 76638
rect 2494 76690 2546 76702
rect 2494 76626 2546 76638
rect 2942 76690 2994 76702
rect 2942 76626 2994 76638
rect 4734 76690 4786 76702
rect 4734 76626 4786 76638
rect 5854 76690 5906 76702
rect 37550 76690 37602 76702
rect 9986 76638 9998 76690
rect 10050 76638 10062 76690
rect 5854 76626 5906 76638
rect 37550 76626 37602 76638
rect 39902 76690 39954 76702
rect 39902 76626 39954 76638
rect 40910 76690 40962 76702
rect 40910 76626 40962 76638
rect 41918 76690 41970 76702
rect 41918 76626 41970 76638
rect 59950 76690 60002 76702
rect 59950 76626 60002 76638
rect 63870 76690 63922 76702
rect 63870 76626 63922 76638
rect 67790 76690 67842 76702
rect 67790 76626 67842 76638
rect 72494 76690 72546 76702
rect 72494 76626 72546 76638
rect 3502 76578 3554 76590
rect 31726 76578 31778 76590
rect 7522 76526 7534 76578
rect 7586 76526 7598 76578
rect 12338 76526 12350 76578
rect 12402 76526 12414 76578
rect 23538 76526 23550 76578
rect 23602 76526 23614 76578
rect 27458 76526 27470 76578
rect 27522 76526 27534 76578
rect 30594 76526 30606 76578
rect 30658 76526 30670 76578
rect 3502 76514 3554 76526
rect 31726 76514 31778 76526
rect 31838 76578 31890 76590
rect 35982 76578 36034 76590
rect 48750 76578 48802 76590
rect 52670 76578 52722 76590
rect 34626 76526 34638 76578
rect 34690 76526 34702 76578
rect 38994 76526 39006 76578
rect 39058 76526 39070 76578
rect 43362 76526 43374 76578
rect 43426 76526 43438 76578
rect 47618 76526 47630 76578
rect 47682 76526 47694 76578
rect 51538 76526 51550 76578
rect 51602 76526 51614 76578
rect 61618 76526 61630 76578
rect 61682 76526 61694 76578
rect 65538 76526 65550 76578
rect 65602 76526 65614 76578
rect 69570 76526 69582 76578
rect 69634 76526 69646 76578
rect 73938 76526 73950 76578
rect 74002 76526 74014 76578
rect 31838 76514 31890 76526
rect 35982 76514 36034 76526
rect 48750 76514 48802 76526
rect 52670 76514 52722 76526
rect 3614 76466 3666 76478
rect 3614 76402 3666 76414
rect 4398 76466 4450 76478
rect 4398 76402 4450 76414
rect 4734 76466 4786 76478
rect 6638 76466 6690 76478
rect 6290 76414 6302 76466
rect 6354 76414 6366 76466
rect 4734 76402 4786 76414
rect 6638 76402 6690 76414
rect 6862 76466 6914 76478
rect 6862 76402 6914 76414
rect 10446 76466 10498 76478
rect 10446 76402 10498 76414
rect 10558 76466 10610 76478
rect 10558 76402 10610 76414
rect 10670 76466 10722 76478
rect 16706 76414 16718 76466
rect 16770 76414 16782 76466
rect 17714 76414 17726 76466
rect 17778 76414 17790 76466
rect 24322 76414 24334 76466
rect 24386 76414 24398 76466
rect 28130 76414 28142 76466
rect 28194 76414 28206 76466
rect 32050 76414 32062 76466
rect 32114 76414 32126 76466
rect 10670 76402 10722 76414
rect 6750 76354 6802 76366
rect 33182 76354 33234 76366
rect 35646 76354 35698 76366
rect 8866 76302 8878 76354
rect 8930 76302 8942 76354
rect 11554 76302 11566 76354
rect 11618 76302 11630 76354
rect 13794 76302 13806 76354
rect 13858 76302 13870 76354
rect 15922 76302 15934 76354
rect 15986 76302 15998 76354
rect 18498 76302 18510 76354
rect 18562 76302 18574 76354
rect 20626 76302 20638 76354
rect 20690 76302 20702 76354
rect 21410 76302 21422 76354
rect 21474 76302 21486 76354
rect 25330 76302 25342 76354
rect 25394 76302 25406 76354
rect 29474 76302 29486 76354
rect 29538 76302 29550 76354
rect 33618 76302 33630 76354
rect 33682 76302 33694 76354
rect 6750 76290 6802 76302
rect 33182 76290 33234 76302
rect 35646 76290 35698 76302
rect 37102 76354 37154 76366
rect 41358 76354 41410 76366
rect 37986 76302 37998 76354
rect 38050 76302 38062 76354
rect 42354 76302 42366 76354
rect 42418 76302 42430 76354
rect 46610 76302 46622 76354
rect 46674 76302 46686 76354
rect 50530 76302 50542 76354
rect 50594 76302 50606 76354
rect 60610 76302 60622 76354
rect 60674 76302 60686 76354
rect 64530 76302 64542 76354
rect 64594 76302 64606 76354
rect 68562 76302 68574 76354
rect 68626 76302 68638 76354
rect 72930 76302 72942 76354
rect 72994 76302 73006 76354
rect 37102 76290 37154 76302
rect 41358 76290 41410 76302
rect 3726 76242 3778 76254
rect 3726 76178 3778 76190
rect 4622 76242 4674 76254
rect 31266 76190 31278 76242
rect 31330 76190 31342 76242
rect 4622 76178 4674 76190
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 2046 75906 2098 75918
rect 37314 75854 37326 75906
rect 37378 75903 37390 75906
rect 37986 75903 37998 75906
rect 37378 75857 37998 75903
rect 37378 75854 37390 75857
rect 37986 75854 37998 75857
rect 38050 75854 38062 75906
rect 2046 75842 2098 75854
rect 3614 75794 3666 75806
rect 29822 75794 29874 75806
rect 36542 75794 36594 75806
rect 3614 75730 3666 75742
rect 4062 75738 4114 75750
rect 6066 75742 6078 75794
rect 6130 75742 6142 75794
rect 8194 75742 8206 75794
rect 8258 75742 8270 75794
rect 12898 75742 12910 75794
rect 12962 75742 12974 75794
rect 14578 75742 14590 75794
rect 14642 75742 14654 75794
rect 16818 75742 16830 75794
rect 16882 75742 16894 75794
rect 19394 75742 19406 75794
rect 19458 75742 19470 75794
rect 22978 75742 22990 75794
rect 23042 75742 23054 75794
rect 25106 75742 25118 75794
rect 25170 75742 25182 75794
rect 28018 75742 28030 75794
rect 28082 75742 28094 75794
rect 31042 75742 31054 75794
rect 31106 75742 31118 75794
rect 29822 75730 29874 75742
rect 36542 75730 36594 75742
rect 38334 75794 38386 75806
rect 38334 75730 38386 75742
rect 38782 75794 38834 75806
rect 38782 75730 38834 75742
rect 40126 75794 40178 75806
rect 40126 75730 40178 75742
rect 55022 75794 55074 75806
rect 77198 75794 77250 75806
rect 55458 75742 55470 75794
rect 55522 75742 55534 75794
rect 74946 75742 74958 75794
rect 75010 75742 75022 75794
rect 55022 75730 55074 75742
rect 77198 75730 77250 75742
rect 4062 75674 4114 75686
rect 4286 75682 4338 75694
rect 4286 75618 4338 75630
rect 4510 75682 4562 75694
rect 13582 75682 13634 75694
rect 21758 75682 21810 75694
rect 31950 75682 32002 75694
rect 8978 75630 8990 75682
rect 9042 75630 9054 75682
rect 10098 75630 10110 75682
rect 10162 75630 10174 75682
rect 17490 75630 17502 75682
rect 17554 75630 17566 75682
rect 22306 75630 22318 75682
rect 22370 75630 22382 75682
rect 28690 75630 28702 75682
rect 28754 75630 28766 75682
rect 30930 75630 30942 75682
rect 30994 75630 31006 75682
rect 32386 75630 32398 75682
rect 32450 75630 32462 75682
rect 32834 75630 32846 75682
rect 32898 75630 32910 75682
rect 34178 75630 34190 75682
rect 34242 75630 34254 75682
rect 34962 75630 34974 75682
rect 35026 75630 35038 75682
rect 4510 75618 4562 75630
rect 13582 75618 13634 75630
rect 21758 75618 21810 75630
rect 31950 75618 32002 75630
rect 4958 75570 5010 75582
rect 13918 75570 13970 75582
rect 4722 75518 4734 75570
rect 4786 75518 4798 75570
rect 10770 75518 10782 75570
rect 10834 75518 10846 75570
rect 4958 75506 5010 75518
rect 13918 75506 13970 75518
rect 18622 75570 18674 75582
rect 31390 75570 31442 75582
rect 33406 75570 33458 75582
rect 20402 75518 20414 75570
rect 20466 75518 20478 75570
rect 32946 75518 32958 75570
rect 33010 75518 33022 75570
rect 18622 75506 18674 75518
rect 31390 75506 31442 75518
rect 33406 75506 33458 75518
rect 36094 75570 36146 75582
rect 56466 75518 56478 75570
rect 56530 75518 56542 75570
rect 76290 75518 76302 75570
rect 76354 75518 76366 75570
rect 36094 75506 36146 75518
rect 2830 75458 2882 75470
rect 2830 75394 2882 75406
rect 4510 75458 4562 75470
rect 4510 75394 4562 75406
rect 9550 75458 9602 75470
rect 9550 75394 9602 75406
rect 13806 75458 13858 75470
rect 13806 75394 13858 75406
rect 18174 75458 18226 75470
rect 18174 75394 18226 75406
rect 18286 75458 18338 75470
rect 18286 75394 18338 75406
rect 18398 75458 18450 75470
rect 35758 75458 35810 75470
rect 25778 75406 25790 75458
rect 25842 75406 25854 75458
rect 18398 75394 18450 75406
rect 35758 75394 35810 75406
rect 37438 75458 37490 75470
rect 37438 75394 37490 75406
rect 37886 75458 37938 75470
rect 37886 75394 37938 75406
rect 39230 75458 39282 75470
rect 39230 75394 39282 75406
rect 39678 75458 39730 75470
rect 39678 75394 39730 75406
rect 40574 75458 40626 75470
rect 40574 75394 40626 75406
rect 41022 75458 41074 75470
rect 41022 75394 41074 75406
rect 41470 75458 41522 75470
rect 41470 75394 41522 75406
rect 41918 75458 41970 75470
rect 41918 75394 41970 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 2382 75122 2434 75134
rect 2382 75058 2434 75070
rect 12350 75122 12402 75134
rect 12350 75058 12402 75070
rect 35422 75122 35474 75134
rect 35422 75058 35474 75070
rect 35870 75122 35922 75134
rect 35870 75058 35922 75070
rect 38558 75122 38610 75134
rect 38558 75058 38610 75070
rect 39454 75122 39506 75134
rect 39454 75058 39506 75070
rect 7758 75010 7810 75022
rect 7758 74946 7810 74958
rect 11342 75010 11394 75022
rect 11342 74946 11394 74958
rect 13022 75010 13074 75022
rect 13022 74946 13074 74958
rect 13134 75010 13186 75022
rect 24894 75010 24946 75022
rect 33742 75010 33794 75022
rect 18722 74958 18734 75010
rect 18786 74958 18798 75010
rect 27794 74958 27806 75010
rect 27858 74958 27870 75010
rect 31826 74958 31838 75010
rect 31890 74958 31902 75010
rect 13134 74946 13186 74958
rect 24894 74946 24946 74958
rect 33742 74946 33794 74958
rect 8430 74898 8482 74910
rect 3154 74846 3166 74898
rect 3218 74846 3230 74898
rect 6850 74846 6862 74898
rect 6914 74846 6926 74898
rect 8430 74834 8482 74846
rect 8766 74898 8818 74910
rect 8766 74834 8818 74846
rect 8990 74898 9042 74910
rect 11454 74898 11506 74910
rect 11106 74846 11118 74898
rect 11170 74846 11182 74898
rect 8990 74834 9042 74846
rect 11454 74834 11506 74846
rect 12574 74898 12626 74910
rect 24222 74898 24274 74910
rect 16930 74846 16942 74898
rect 16994 74846 17006 74898
rect 20290 74846 20302 74898
rect 20354 74846 20366 74898
rect 12574 74834 12626 74846
rect 24222 74834 24274 74846
rect 24446 74898 24498 74910
rect 24446 74834 24498 74846
rect 24670 74898 24722 74910
rect 31166 74898 31218 74910
rect 34302 74898 34354 74910
rect 28578 74846 28590 74898
rect 28642 74846 28654 74898
rect 29698 74846 29710 74898
rect 29762 74846 29774 74898
rect 30818 74846 30830 74898
rect 30882 74846 30894 74898
rect 31938 74846 31950 74898
rect 32002 74846 32014 74898
rect 32386 74846 32398 74898
rect 32450 74846 32462 74898
rect 34514 74846 34526 74898
rect 34578 74846 34590 74898
rect 24670 74834 24722 74846
rect 31166 74834 31218 74846
rect 34302 74834 34354 74846
rect 1934 74786 1986 74798
rect 8542 74786 8594 74798
rect 3826 74734 3838 74786
rect 3890 74734 3902 74786
rect 6066 74734 6078 74786
rect 6130 74734 6142 74786
rect 1934 74722 1986 74734
rect 8542 74722 8594 74734
rect 10558 74786 10610 74798
rect 10558 74722 10610 74734
rect 13358 74786 13410 74798
rect 19854 74786 19906 74798
rect 23214 74786 23266 74798
rect 29038 74786 29090 74798
rect 14018 74734 14030 74786
rect 14082 74734 14094 74786
rect 16146 74734 16158 74786
rect 16210 74734 16222 74786
rect 17714 74734 17726 74786
rect 17778 74734 17790 74786
rect 21074 74734 21086 74786
rect 21138 74734 21150 74786
rect 25666 74734 25678 74786
rect 25730 74734 25742 74786
rect 13358 74722 13410 74734
rect 19854 74722 19906 74734
rect 23214 74722 23266 74734
rect 29038 74722 29090 74734
rect 32846 74786 32898 74798
rect 32846 74722 32898 74734
rect 34974 74786 35026 74798
rect 34974 74722 35026 74734
rect 36318 74786 36370 74798
rect 36318 74722 36370 74734
rect 36766 74786 36818 74798
rect 36766 74722 36818 74734
rect 37214 74786 37266 74798
rect 37214 74722 37266 74734
rect 37662 74786 37714 74798
rect 37662 74722 37714 74734
rect 38110 74786 38162 74798
rect 38110 74722 38162 74734
rect 39006 74786 39058 74798
rect 39006 74722 39058 74734
rect 39902 74786 39954 74798
rect 39902 74722 39954 74734
rect 40350 74786 40402 74798
rect 40350 74722 40402 74734
rect 40798 74786 40850 74798
rect 40798 74722 40850 74734
rect 41470 74786 41522 74798
rect 41470 74722 41522 74734
rect 2830 74674 2882 74686
rect 2830 74610 2882 74622
rect 3166 74674 3218 74686
rect 3166 74610 3218 74622
rect 7534 74674 7586 74686
rect 7534 74610 7586 74622
rect 7870 74674 7922 74686
rect 10334 74674 10386 74686
rect 24782 74674 24834 74686
rect 9986 74622 9998 74674
rect 10050 74622 10062 74674
rect 11890 74622 11902 74674
rect 11954 74622 11966 74674
rect 7870 74610 7922 74622
rect 10334 74610 10386 74622
rect 24782 74610 24834 74622
rect 33854 74674 33906 74686
rect 33854 74610 33906 74622
rect 34078 74674 34130 74686
rect 37538 74622 37550 74674
rect 37602 74671 37614 74674
rect 38994 74671 39006 74674
rect 37602 74625 39006 74671
rect 37602 74622 37614 74625
rect 38994 74622 39006 74625
rect 39058 74622 39070 74674
rect 34078 74610 34130 74622
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 7086 74338 7138 74350
rect 2930 74286 2942 74338
rect 2994 74335 3006 74338
rect 3266 74335 3278 74338
rect 2994 74289 3278 74335
rect 2994 74286 3006 74289
rect 3266 74286 3278 74289
rect 3330 74286 3342 74338
rect 7086 74274 7138 74286
rect 9662 74338 9714 74350
rect 11790 74338 11842 74350
rect 11218 74286 11230 74338
rect 11282 74286 11294 74338
rect 37314 74286 37326 74338
rect 37378 74335 37390 74338
rect 38098 74335 38110 74338
rect 37378 74289 38110 74335
rect 37378 74286 37390 74289
rect 38098 74286 38110 74289
rect 38162 74286 38174 74338
rect 38658 74286 38670 74338
rect 38722 74335 38734 74338
rect 39890 74335 39902 74338
rect 38722 74289 39902 74335
rect 38722 74286 38734 74289
rect 39890 74286 39902 74289
rect 39954 74286 39966 74338
rect 9662 74274 9714 74286
rect 11790 74274 11842 74286
rect 2158 74226 2210 74238
rect 2158 74162 2210 74174
rect 2606 74226 2658 74238
rect 2606 74162 2658 74174
rect 3054 74226 3106 74238
rect 3054 74162 3106 74174
rect 4846 74226 4898 74238
rect 31390 74226 31442 74238
rect 5954 74174 5966 74226
rect 6018 74174 6030 74226
rect 14466 74174 14478 74226
rect 14530 74174 14542 74226
rect 16594 74174 16606 74226
rect 16658 74174 16670 74226
rect 17938 74174 17950 74226
rect 18002 74174 18014 74226
rect 20066 74174 20078 74226
rect 20130 74174 20142 74226
rect 26338 74174 26350 74226
rect 26402 74174 26414 74226
rect 27010 74174 27022 74226
rect 27074 74174 27086 74226
rect 30594 74174 30606 74226
rect 30658 74174 30670 74226
rect 4846 74162 4898 74174
rect 31390 74162 31442 74174
rect 32174 74226 32226 74238
rect 32174 74162 32226 74174
rect 36766 74226 36818 74238
rect 36766 74162 36818 74174
rect 37886 74226 37938 74238
rect 37886 74162 37938 74174
rect 38334 74226 38386 74238
rect 38334 74162 38386 74174
rect 38782 74226 38834 74238
rect 38782 74162 38834 74174
rect 4734 74114 4786 74126
rect 4386 74062 4398 74114
rect 4450 74062 4462 74114
rect 4734 74050 4786 74062
rect 4958 74114 5010 74126
rect 4958 74050 5010 74062
rect 6974 74114 7026 74126
rect 7758 74114 7810 74126
rect 8878 74114 8930 74126
rect 7634 74062 7646 74114
rect 7698 74062 7710 74114
rect 7970 74062 7982 74114
rect 8034 74062 8046 74114
rect 8642 74062 8654 74114
rect 8706 74062 8718 74114
rect 6974 74050 7026 74062
rect 7758 74050 7810 74062
rect 8878 74050 8930 74062
rect 9774 74114 9826 74126
rect 9774 74050 9826 74062
rect 9998 74114 10050 74126
rect 11006 74114 11058 74126
rect 10658 74062 10670 74114
rect 10722 74062 10734 74114
rect 9998 74050 10050 74062
rect 11006 74050 11058 74062
rect 11118 74114 11170 74126
rect 11118 74050 11170 74062
rect 11342 74114 11394 74126
rect 11342 74050 11394 74062
rect 12014 74114 12066 74126
rect 22094 74114 22146 74126
rect 33630 74114 33682 74126
rect 35982 74114 36034 74126
rect 13794 74062 13806 74114
rect 13858 74062 13870 74114
rect 17154 74062 17166 74114
rect 17218 74062 17230 74114
rect 23426 74062 23438 74114
rect 23490 74062 23502 74114
rect 30258 74062 30270 74114
rect 30322 74062 30334 74114
rect 32498 74062 32510 74114
rect 32562 74062 32574 74114
rect 32946 74062 32958 74114
rect 33010 74062 33022 74114
rect 34402 74062 34414 74114
rect 34466 74062 34478 74114
rect 35186 74062 35198 74114
rect 35250 74062 35262 74114
rect 12014 74050 12066 74062
rect 22094 74050 22146 74062
rect 33630 74050 33682 74062
rect 35982 74050 36034 74062
rect 3502 74002 3554 74014
rect 3502 73938 3554 73950
rect 3950 74002 4002 74014
rect 3950 73938 4002 73950
rect 7422 74002 7474 74014
rect 7422 73938 7474 73950
rect 8990 74002 9042 74014
rect 8990 73938 9042 73950
rect 10110 74002 10162 74014
rect 10110 73938 10162 73950
rect 12686 74002 12738 74014
rect 12686 73938 12738 73950
rect 12798 74002 12850 74014
rect 12798 73938 12850 73950
rect 12910 74002 12962 74014
rect 12910 73938 12962 73950
rect 20862 74002 20914 74014
rect 20862 73938 20914 73950
rect 21646 74002 21698 74014
rect 21646 73938 21698 73950
rect 22318 74002 22370 74014
rect 22318 73938 22370 73950
rect 22766 74002 22818 74014
rect 30942 74002 30994 74014
rect 24098 73950 24110 74002
rect 24162 73950 24174 74002
rect 28354 73950 28366 74002
rect 28418 73950 28430 74002
rect 22766 73938 22818 73950
rect 30942 73938 30994 73950
rect 37438 74002 37490 74014
rect 37438 73938 37490 73950
rect 6414 73890 6466 73902
rect 6414 73826 6466 73838
rect 20526 73890 20578 73902
rect 20526 73826 20578 73838
rect 20750 73890 20802 73902
rect 20750 73826 20802 73838
rect 21870 73890 21922 73902
rect 21870 73826 21922 73838
rect 22430 73890 22482 73902
rect 36318 73890 36370 73902
rect 33170 73838 33182 73890
rect 33234 73838 33246 73890
rect 22430 73826 22482 73838
rect 36318 73826 36370 73838
rect 39230 73890 39282 73902
rect 39230 73826 39282 73838
rect 39678 73890 39730 73902
rect 39678 73826 39730 73838
rect 40126 73890 40178 73902
rect 40126 73826 40178 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 1934 73554 1986 73566
rect 1934 73490 1986 73502
rect 2382 73554 2434 73566
rect 2382 73490 2434 73502
rect 7646 73554 7698 73566
rect 7646 73490 7698 73502
rect 23998 73554 24050 73566
rect 23998 73490 24050 73502
rect 35534 73554 35586 73566
rect 35534 73490 35586 73502
rect 36430 73554 36482 73566
rect 36430 73490 36482 73502
rect 37326 73554 37378 73566
rect 37326 73490 37378 73502
rect 4174 73442 4226 73454
rect 4174 73378 4226 73390
rect 6750 73442 6802 73454
rect 6750 73378 6802 73390
rect 8990 73442 9042 73454
rect 18510 73442 18562 73454
rect 10210 73390 10222 73442
rect 10274 73390 10286 73442
rect 14802 73390 14814 73442
rect 14866 73390 14878 73442
rect 8990 73378 9042 73390
rect 18510 73378 18562 73390
rect 19182 73442 19234 73454
rect 19182 73378 19234 73390
rect 29150 73442 29202 73454
rect 29150 73378 29202 73390
rect 30494 73442 30546 73454
rect 30494 73378 30546 73390
rect 32398 73442 32450 73454
rect 32398 73378 32450 73390
rect 36878 73442 36930 73454
rect 36878 73378 36930 73390
rect 5182 73330 5234 73342
rect 4498 73278 4510 73330
rect 4562 73278 4574 73330
rect 5182 73266 5234 73278
rect 5406 73330 5458 73342
rect 5406 73266 5458 73278
rect 6190 73330 6242 73342
rect 6190 73266 6242 73278
rect 6414 73330 6466 73342
rect 6414 73266 6466 73278
rect 7198 73330 7250 73342
rect 7198 73266 7250 73278
rect 7870 73330 7922 73342
rect 7870 73266 7922 73278
rect 8878 73330 8930 73342
rect 17950 73330 18002 73342
rect 10658 73278 10670 73330
rect 10722 73278 10734 73330
rect 11330 73278 11342 73330
rect 11394 73278 11406 73330
rect 13010 73278 13022 73330
rect 13074 73278 13086 73330
rect 14018 73278 14030 73330
rect 14082 73278 14094 73330
rect 17714 73278 17726 73330
rect 17778 73278 17790 73330
rect 8878 73266 8930 73278
rect 17950 73266 18002 73278
rect 18174 73330 18226 73342
rect 23662 73330 23714 73342
rect 19394 73278 19406 73330
rect 19458 73278 19470 73330
rect 20178 73278 20190 73330
rect 20242 73278 20254 73330
rect 18174 73266 18226 73278
rect 23662 73266 23714 73278
rect 23998 73330 24050 73342
rect 23998 73266 24050 73278
rect 24334 73330 24386 73342
rect 29374 73330 29426 73342
rect 28578 73278 28590 73330
rect 28642 73278 28654 73330
rect 24334 73266 24386 73278
rect 29374 73266 29426 73278
rect 29710 73330 29762 73342
rect 29710 73266 29762 73278
rect 29822 73330 29874 73342
rect 31490 73278 31502 73330
rect 31554 73278 31566 73330
rect 33954 73278 33966 73330
rect 34018 73278 34030 73330
rect 29822 73266 29874 73278
rect 2830 73218 2882 73230
rect 2830 73154 2882 73166
rect 3278 73218 3330 73230
rect 3278 73154 3330 73166
rect 3726 73218 3778 73230
rect 3726 73154 3778 73166
rect 4286 73218 4338 73230
rect 4286 73154 4338 73166
rect 6638 73218 6690 73230
rect 6638 73154 6690 73166
rect 7758 73218 7810 73230
rect 22990 73218 23042 73230
rect 11778 73166 11790 73218
rect 11842 73166 11854 73218
rect 12786 73166 12798 73218
rect 12850 73166 12862 73218
rect 16930 73166 16942 73218
rect 16994 73166 17006 73218
rect 20850 73166 20862 73218
rect 20914 73166 20926 73218
rect 7758 73154 7810 73166
rect 22990 73154 23042 73166
rect 24894 73218 24946 73230
rect 32846 73218 32898 73230
rect 34638 73218 34690 73230
rect 25666 73166 25678 73218
rect 25730 73166 25742 73218
rect 27794 73166 27806 73218
rect 27858 73166 27870 73218
rect 31714 73166 31726 73218
rect 31778 73166 31790 73218
rect 33730 73166 33742 73218
rect 33794 73166 33806 73218
rect 24894 73154 24946 73166
rect 32846 73154 32898 73166
rect 34638 73154 34690 73166
rect 35086 73218 35138 73230
rect 35086 73154 35138 73166
rect 35982 73218 36034 73230
rect 35982 73154 36034 73166
rect 37774 73218 37826 73230
rect 37774 73154 37826 73166
rect 38222 73218 38274 73230
rect 38222 73154 38274 73166
rect 38670 73218 38722 73230
rect 38670 73154 38722 73166
rect 39118 73218 39170 73230
rect 39118 73154 39170 73166
rect 39566 73218 39618 73230
rect 39566 73154 39618 73166
rect 5070 73106 5122 73118
rect 5070 73042 5122 73054
rect 5518 73106 5570 73118
rect 5518 73042 5570 73054
rect 8542 73106 8594 73118
rect 8542 73042 8594 73054
rect 8654 73106 8706 73118
rect 8654 73042 8706 73054
rect 10222 73106 10274 73118
rect 18398 73106 18450 73118
rect 30270 73106 30322 73118
rect 13346 73054 13358 73106
rect 13410 73054 13422 73106
rect 29138 73054 29150 73106
rect 29202 73054 29214 73106
rect 35522 73054 35534 73106
rect 35586 73103 35598 73106
rect 35970 73103 35982 73106
rect 35586 73057 35982 73103
rect 35586 73054 35598 73057
rect 35970 73054 35982 73057
rect 36034 73054 36046 73106
rect 10222 73042 10274 73054
rect 18398 73042 18450 73054
rect 30270 73042 30322 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 6302 72770 6354 72782
rect 3378 72718 3390 72770
rect 3442 72767 3454 72770
rect 3826 72767 3838 72770
rect 3442 72721 3838 72767
rect 3442 72718 3454 72721
rect 3826 72718 3838 72721
rect 3890 72767 3902 72770
rect 4498 72767 4510 72770
rect 3890 72721 4510 72767
rect 3890 72718 3902 72721
rect 4498 72718 4510 72721
rect 4562 72718 4574 72770
rect 6302 72706 6354 72718
rect 7086 72770 7138 72782
rect 19742 72770 19794 72782
rect 7410 72718 7422 72770
rect 7474 72718 7486 72770
rect 7086 72706 7138 72718
rect 19742 72706 19794 72718
rect 30270 72770 30322 72782
rect 33954 72718 33966 72770
rect 34018 72767 34030 72770
rect 34626 72767 34638 72770
rect 34018 72721 34638 72767
rect 34018 72718 34030 72721
rect 34626 72718 34638 72721
rect 34690 72767 34702 72770
rect 34962 72767 34974 72770
rect 34690 72721 34974 72767
rect 34690 72718 34702 72721
rect 34962 72718 34974 72721
rect 35026 72718 35038 72770
rect 30270 72706 30322 72718
rect 2046 72658 2098 72670
rect 2046 72594 2098 72606
rect 2942 72658 2994 72670
rect 2942 72594 2994 72606
rect 3390 72658 3442 72670
rect 3390 72594 3442 72606
rect 4286 72658 4338 72670
rect 11678 72658 11730 72670
rect 20414 72658 20466 72670
rect 25118 72658 25170 72670
rect 30494 72658 30546 72670
rect 9986 72606 9998 72658
rect 10050 72606 10062 72658
rect 12002 72606 12014 72658
rect 12066 72606 12078 72658
rect 21634 72606 21646 72658
rect 21698 72606 21710 72658
rect 23762 72606 23774 72658
rect 23826 72606 23838 72658
rect 28018 72606 28030 72658
rect 28082 72606 28094 72658
rect 4286 72594 4338 72606
rect 11678 72594 11730 72606
rect 20414 72594 20466 72606
rect 25118 72594 25170 72606
rect 30494 72594 30546 72606
rect 32062 72658 32114 72670
rect 32062 72594 32114 72606
rect 34638 72658 34690 72670
rect 34638 72594 34690 72606
rect 35646 72658 35698 72670
rect 35646 72594 35698 72606
rect 36430 72658 36482 72670
rect 36430 72594 36482 72606
rect 37886 72658 37938 72670
rect 37886 72594 37938 72606
rect 3838 72546 3890 72558
rect 3838 72482 3890 72494
rect 6862 72546 6914 72558
rect 6862 72482 6914 72494
rect 7982 72546 8034 72558
rect 7982 72482 8034 72494
rect 8206 72546 8258 72558
rect 18286 72546 18338 72558
rect 9090 72494 9102 72546
rect 9154 72494 9166 72546
rect 12226 72494 12238 72546
rect 12290 72494 12302 72546
rect 17378 72494 17390 72546
rect 17442 72494 17454 72546
rect 8206 72482 8258 72494
rect 18286 72482 18338 72494
rect 18510 72546 18562 72558
rect 18510 72482 18562 72494
rect 20302 72546 20354 72558
rect 30718 72546 30770 72558
rect 24434 72494 24446 72546
rect 24498 72494 24510 72546
rect 28802 72494 28814 72546
rect 28866 72494 28878 72546
rect 20302 72482 20354 72494
rect 30718 72482 30770 72494
rect 30830 72546 30882 72558
rect 30830 72482 30882 72494
rect 31838 72546 31890 72558
rect 31838 72482 31890 72494
rect 32622 72546 32674 72558
rect 32622 72482 32674 72494
rect 33518 72546 33570 72558
rect 33518 72482 33570 72494
rect 38334 72546 38386 72558
rect 38334 72482 38386 72494
rect 38782 72546 38834 72558
rect 38782 72482 38834 72494
rect 4734 72434 4786 72446
rect 4734 72370 4786 72382
rect 5966 72434 6018 72446
rect 5966 72370 6018 72382
rect 11006 72434 11058 72446
rect 11006 72370 11058 72382
rect 11118 72434 11170 72446
rect 11118 72370 11170 72382
rect 13694 72434 13746 72446
rect 18062 72434 18114 72446
rect 16706 72382 16718 72434
rect 16770 72382 16782 72434
rect 13694 72370 13746 72382
rect 18062 72370 18114 72382
rect 20638 72434 20690 72446
rect 20638 72370 20690 72382
rect 20862 72434 20914 72446
rect 20862 72370 20914 72382
rect 32958 72434 33010 72446
rect 32958 72370 33010 72382
rect 35982 72434 36034 72446
rect 35982 72370 36034 72382
rect 2494 72322 2546 72334
rect 2494 72258 2546 72270
rect 4846 72322 4898 72334
rect 4846 72258 4898 72270
rect 5070 72322 5122 72334
rect 5070 72258 5122 72270
rect 6190 72322 6242 72334
rect 10782 72322 10834 72334
rect 8530 72270 8542 72322
rect 8594 72270 8606 72322
rect 6190 72258 6242 72270
rect 10782 72258 10834 72270
rect 13806 72322 13858 72334
rect 18398 72322 18450 72334
rect 14466 72270 14478 72322
rect 14530 72270 14542 72322
rect 13806 72258 13858 72270
rect 18398 72258 18450 72270
rect 18622 72322 18674 72334
rect 18622 72258 18674 72270
rect 19518 72322 19570 72334
rect 19518 72258 19570 72270
rect 19630 72322 19682 72334
rect 29598 72322 29650 72334
rect 25778 72270 25790 72322
rect 25842 72270 25854 72322
rect 19630 72258 19682 72270
rect 29598 72258 29650 72270
rect 30382 72322 30434 72334
rect 33630 72322 33682 72334
rect 31490 72270 31502 72322
rect 31554 72270 31566 72322
rect 30382 72258 30434 72270
rect 33630 72258 33682 72270
rect 33854 72322 33906 72334
rect 33854 72258 33906 72270
rect 34190 72322 34242 72334
rect 34190 72258 34242 72270
rect 35086 72322 35138 72334
rect 35086 72258 35138 72270
rect 37438 72322 37490 72334
rect 37438 72258 37490 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 1934 71986 1986 71998
rect 1934 71922 1986 71934
rect 2382 71986 2434 71998
rect 2382 71922 2434 71934
rect 5630 71986 5682 71998
rect 5630 71922 5682 71934
rect 9774 71986 9826 71998
rect 9774 71922 9826 71934
rect 18062 71986 18114 71998
rect 18062 71922 18114 71934
rect 18286 71986 18338 71998
rect 18286 71922 18338 71934
rect 27246 71986 27298 71998
rect 27246 71922 27298 71934
rect 32398 71986 32450 71998
rect 32398 71922 32450 71934
rect 34078 71986 34130 71998
rect 34078 71922 34130 71934
rect 36878 71986 36930 71998
rect 36878 71922 36930 71934
rect 37326 71986 37378 71998
rect 37326 71922 37378 71934
rect 5406 71874 5458 71886
rect 5406 71810 5458 71822
rect 5742 71874 5794 71886
rect 5742 71810 5794 71822
rect 6526 71874 6578 71886
rect 33854 71874 33906 71886
rect 8082 71822 8094 71874
rect 8146 71822 8158 71874
rect 29362 71822 29374 71874
rect 29426 71822 29438 71874
rect 6526 71810 6578 71822
rect 33854 71810 33906 71822
rect 35086 71874 35138 71886
rect 35086 71810 35138 71822
rect 35534 71874 35586 71886
rect 35534 71810 35586 71822
rect 3390 71762 3442 71774
rect 5966 71762 6018 71774
rect 10670 71762 10722 71774
rect 3826 71710 3838 71762
rect 3890 71710 3902 71762
rect 7186 71710 7198 71762
rect 7250 71710 7262 71762
rect 3390 71698 3442 71710
rect 5966 71698 6018 71710
rect 10670 71698 10722 71710
rect 10782 71762 10834 71774
rect 10782 71698 10834 71710
rect 10894 71762 10946 71774
rect 18734 71762 18786 71774
rect 24894 71762 24946 71774
rect 16706 71710 16718 71762
rect 16770 71710 16782 71762
rect 19170 71710 19182 71762
rect 19234 71710 19246 71762
rect 10894 71698 10946 71710
rect 18734 71698 18786 71710
rect 24894 71698 24946 71710
rect 25678 71762 25730 71774
rect 25678 71698 25730 71710
rect 25902 71762 25954 71774
rect 25902 71698 25954 71710
rect 26350 71762 26402 71774
rect 27582 71762 27634 71774
rect 27458 71710 27470 71762
rect 27522 71710 27534 71762
rect 26350 71698 26402 71710
rect 27582 71698 27634 71710
rect 27694 71762 27746 71774
rect 30046 71762 30098 71774
rect 32286 71762 32338 71774
rect 28690 71710 28702 71762
rect 28754 71710 28766 71762
rect 29138 71710 29150 71762
rect 29202 71710 29214 71762
rect 30594 71710 30606 71762
rect 30658 71710 30670 71762
rect 31378 71710 31390 71762
rect 31442 71710 31454 71762
rect 27694 71698 27746 71710
rect 30046 71698 30098 71710
rect 32286 71698 32338 71710
rect 32622 71762 32674 71774
rect 32622 71698 32674 71710
rect 32846 71762 32898 71774
rect 32846 71698 32898 71710
rect 34190 71762 34242 71774
rect 34190 71698 34242 71710
rect 37774 71762 37826 71774
rect 37774 71698 37826 71710
rect 2830 71650 2882 71662
rect 2830 71586 2882 71598
rect 4286 71650 4338 71662
rect 4286 71586 4338 71598
rect 4846 71650 4898 71662
rect 4846 71586 4898 71598
rect 8542 71650 8594 71662
rect 18174 71650 18226 71662
rect 25790 71650 25842 71662
rect 13346 71598 13358 71650
rect 13410 71598 13422 71650
rect 24210 71598 24222 71650
rect 24274 71598 24286 71650
rect 8542 71586 8594 71598
rect 18174 71586 18226 71598
rect 25790 71586 25842 71598
rect 28366 71650 28418 71662
rect 28366 71586 28418 71598
rect 34638 71650 34690 71662
rect 34638 71586 34690 71598
rect 35982 71650 36034 71662
rect 35982 71586 36034 71598
rect 36430 71650 36482 71662
rect 36430 71586 36482 71598
rect 38222 71650 38274 71662
rect 38222 71586 38274 71598
rect 26798 71538 26850 71550
rect 10210 71486 10222 71538
rect 10274 71486 10286 71538
rect 26798 71474 26850 71486
rect 26910 71538 26962 71550
rect 36418 71486 36430 71538
rect 36482 71535 36494 71538
rect 36642 71535 36654 71538
rect 36482 71489 36654 71535
rect 36482 71486 36494 71489
rect 36642 71486 36654 71489
rect 36706 71486 36718 71538
rect 37426 71486 37438 71538
rect 37490 71535 37502 71538
rect 38322 71535 38334 71538
rect 37490 71489 38334 71535
rect 37490 71486 37502 71489
rect 38322 71486 38334 71489
rect 38386 71486 38398 71538
rect 26910 71474 26962 71486
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 5630 71202 5682 71214
rect 5630 71138 5682 71150
rect 7310 71202 7362 71214
rect 7310 71138 7362 71150
rect 13918 71202 13970 71214
rect 26126 71202 26178 71214
rect 25218 71150 25230 71202
rect 25282 71150 25294 71202
rect 13918 71138 13970 71150
rect 26126 71138 26178 71150
rect 26238 71202 26290 71214
rect 26238 71138 26290 71150
rect 28590 71202 28642 71214
rect 28590 71138 28642 71150
rect 29598 71202 29650 71214
rect 29598 71138 29650 71150
rect 29710 71202 29762 71214
rect 29710 71138 29762 71150
rect 30158 71202 30210 71214
rect 30158 71138 30210 71150
rect 2158 71090 2210 71102
rect 2158 71026 2210 71038
rect 2606 71090 2658 71102
rect 2606 71026 2658 71038
rect 3502 71090 3554 71102
rect 3502 71026 3554 71038
rect 3950 71090 4002 71102
rect 3950 71026 4002 71038
rect 4622 71090 4674 71102
rect 4622 71026 4674 71038
rect 11902 71090 11954 71102
rect 11902 71026 11954 71038
rect 12798 71090 12850 71102
rect 28702 71090 28754 71102
rect 21634 71038 21646 71090
rect 21698 71038 21710 71090
rect 23762 71038 23774 71090
rect 23826 71038 23838 71090
rect 27122 71038 27134 71090
rect 27186 71038 27198 71090
rect 12798 71026 12850 71038
rect 28702 71026 28754 71038
rect 32062 71090 32114 71102
rect 32062 71026 32114 71038
rect 35198 71090 35250 71102
rect 35198 71026 35250 71038
rect 35534 71090 35586 71102
rect 35534 71026 35586 71038
rect 36430 71090 36482 71102
rect 36430 71026 36482 71038
rect 37438 71090 37490 71102
rect 37438 71026 37490 71038
rect 4398 70978 4450 70990
rect 6302 70978 6354 70990
rect 5954 70926 5966 70978
rect 6018 70926 6030 70978
rect 4398 70914 4450 70926
rect 6302 70914 6354 70926
rect 6414 70978 6466 70990
rect 6414 70914 6466 70926
rect 6526 70978 6578 70990
rect 6526 70914 6578 70926
rect 7422 70978 7474 70990
rect 12686 70978 12738 70990
rect 10994 70926 11006 70978
rect 11058 70926 11070 70978
rect 7422 70914 7474 70926
rect 12686 70914 12738 70926
rect 14142 70978 14194 70990
rect 14142 70914 14194 70926
rect 14366 70978 14418 70990
rect 25566 70978 25618 70990
rect 29934 70978 29986 70990
rect 32958 70978 33010 70990
rect 15250 70926 15262 70978
rect 15314 70926 15326 70978
rect 24546 70926 24558 70978
rect 24610 70926 24622 70978
rect 27570 70926 27582 70978
rect 27634 70926 27646 70978
rect 30370 70926 30382 70978
rect 30434 70926 30446 70978
rect 31490 70926 31502 70978
rect 31554 70926 31566 70978
rect 31826 70926 31838 70978
rect 31890 70926 31902 70978
rect 14366 70914 14418 70926
rect 25566 70914 25618 70926
rect 29934 70914 29986 70926
rect 32958 70914 33010 70926
rect 33406 70978 33458 70990
rect 33406 70914 33458 70926
rect 33742 70978 33794 70990
rect 33742 70914 33794 70926
rect 34638 70978 34690 70990
rect 34638 70914 34690 70926
rect 7310 70866 7362 70878
rect 13694 70866 13746 70878
rect 25118 70866 25170 70878
rect 10322 70814 10334 70866
rect 10386 70814 10398 70866
rect 19170 70814 19182 70866
rect 19234 70814 19246 70866
rect 7310 70802 7362 70814
rect 13694 70802 13746 70814
rect 25118 70802 25170 70814
rect 25454 70866 25506 70878
rect 25454 70802 25506 70814
rect 26462 70866 26514 70878
rect 26462 70802 26514 70814
rect 28030 70866 28082 70878
rect 28030 70802 28082 70814
rect 2942 70754 2994 70766
rect 12462 70754 12514 70766
rect 4946 70702 4958 70754
rect 5010 70702 5022 70754
rect 8082 70702 8094 70754
rect 8146 70702 8158 70754
rect 2942 70690 2994 70702
rect 12462 70690 12514 70702
rect 12910 70754 12962 70766
rect 12910 70690 12962 70702
rect 14814 70754 14866 70766
rect 14814 70690 14866 70702
rect 32622 70754 32674 70766
rect 32622 70690 32674 70702
rect 33630 70754 33682 70766
rect 33630 70690 33682 70702
rect 34190 70754 34242 70766
rect 34190 70690 34242 70702
rect 35982 70754 36034 70766
rect 35982 70690 36034 70702
rect 37886 70754 37938 70766
rect 37886 70690 37938 70702
rect 38334 70754 38386 70766
rect 38334 70690 38386 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 4398 70418 4450 70430
rect 4398 70354 4450 70366
rect 5630 70418 5682 70430
rect 5630 70354 5682 70366
rect 5854 70418 5906 70430
rect 5854 70354 5906 70366
rect 6750 70418 6802 70430
rect 6750 70354 6802 70366
rect 8318 70418 8370 70430
rect 8318 70354 8370 70366
rect 8542 70418 8594 70430
rect 8542 70354 8594 70366
rect 18174 70418 18226 70430
rect 18174 70354 18226 70366
rect 18846 70418 18898 70430
rect 18846 70354 18898 70366
rect 23886 70418 23938 70430
rect 23886 70354 23938 70366
rect 24110 70418 24162 70430
rect 24110 70354 24162 70366
rect 29486 70418 29538 70430
rect 29486 70354 29538 70366
rect 33742 70418 33794 70430
rect 33742 70354 33794 70366
rect 35646 70418 35698 70430
rect 35646 70354 35698 70366
rect 36430 70418 36482 70430
rect 36430 70354 36482 70366
rect 2494 70306 2546 70318
rect 29598 70306 29650 70318
rect 6850 70254 6862 70306
rect 6914 70303 6926 70306
rect 7074 70303 7086 70306
rect 6914 70257 7086 70303
rect 6914 70254 6926 70257
rect 7074 70254 7086 70257
rect 7138 70254 7150 70306
rect 2494 70242 2546 70254
rect 29598 70242 29650 70254
rect 29822 70306 29874 70318
rect 29822 70242 29874 70254
rect 35086 70306 35138 70318
rect 35086 70242 35138 70254
rect 2046 70194 2098 70206
rect 2046 70130 2098 70142
rect 2270 70194 2322 70206
rect 2270 70130 2322 70142
rect 3838 70194 3890 70206
rect 3838 70130 3890 70142
rect 5182 70194 5234 70206
rect 8206 70194 8258 70206
rect 18734 70194 18786 70206
rect 24334 70194 24386 70206
rect 29374 70194 29426 70206
rect 32062 70194 32114 70206
rect 7186 70142 7198 70194
rect 7250 70142 7262 70194
rect 8754 70142 8766 70194
rect 8818 70142 8830 70194
rect 10098 70142 10110 70194
rect 10162 70142 10174 70194
rect 13458 70142 13470 70194
rect 13522 70142 13534 70194
rect 18162 70142 18174 70194
rect 18226 70142 18238 70194
rect 18498 70142 18510 70194
rect 18562 70142 18574 70194
rect 23090 70142 23102 70194
rect 23154 70142 23166 70194
rect 28578 70142 28590 70194
rect 28642 70142 28654 70194
rect 29138 70142 29150 70194
rect 29202 70142 29214 70194
rect 31042 70142 31054 70194
rect 31106 70142 31118 70194
rect 5182 70130 5234 70142
rect 8206 70130 8258 70142
rect 18734 70130 18786 70142
rect 24334 70130 24386 70142
rect 29374 70130 29426 70142
rect 32062 70130 32114 70142
rect 32286 70194 32338 70206
rect 33518 70194 33570 70206
rect 32610 70142 32622 70194
rect 32674 70142 32686 70194
rect 32286 70130 32338 70142
rect 33518 70130 33570 70142
rect 33854 70194 33906 70206
rect 33854 70130 33906 70142
rect 34078 70194 34130 70206
rect 34078 70130 34130 70142
rect 36990 70194 37042 70206
rect 36990 70130 37042 70142
rect 37326 70194 37378 70206
rect 37326 70130 37378 70142
rect 2382 70082 2434 70094
rect 2382 70018 2434 70030
rect 3054 70082 3106 70094
rect 3054 70018 3106 70030
rect 3390 70082 3442 70094
rect 3390 70018 3442 70030
rect 4734 70082 4786 70094
rect 4734 70018 4786 70030
rect 5742 70082 5794 70094
rect 7534 70082 7586 70094
rect 7298 70030 7310 70082
rect 7362 70030 7374 70082
rect 5742 70018 5794 70030
rect 7534 70018 7586 70030
rect 8430 70082 8482 70094
rect 16382 70082 16434 70094
rect 10770 70030 10782 70082
rect 10834 70030 10846 70082
rect 12898 70030 12910 70082
rect 12962 70030 12974 70082
rect 14242 70030 14254 70082
rect 14306 70030 14318 70082
rect 8430 70018 8482 70030
rect 16382 70018 16434 70030
rect 17614 70082 17666 70094
rect 17614 70018 17666 70030
rect 17950 70082 18002 70094
rect 17950 70018 18002 70030
rect 19518 70082 19570 70094
rect 24222 70082 24274 70094
rect 20178 70030 20190 70082
rect 20242 70030 20254 70082
rect 22418 70030 22430 70082
rect 22482 70030 22494 70082
rect 19518 70018 19570 70030
rect 24222 70018 24274 70030
rect 24894 70082 24946 70094
rect 31502 70082 31554 70094
rect 25666 70030 25678 70082
rect 25730 70030 25742 70082
rect 27794 70030 27806 70082
rect 27858 70030 27870 70082
rect 31154 70030 31166 70082
rect 31218 70030 31230 70082
rect 24894 70018 24946 70030
rect 31502 70018 31554 70030
rect 32174 70082 32226 70094
rect 32174 70018 32226 70030
rect 34638 70082 34690 70094
rect 34638 70018 34690 70030
rect 35982 70082 36034 70094
rect 35982 70018 36034 70030
rect 35970 69918 35982 69970
rect 36034 69967 36046 69970
rect 36642 69967 36654 69970
rect 36034 69921 36654 69967
rect 36034 69918 36046 69921
rect 36642 69918 36654 69921
rect 36706 69918 36718 69970
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 5854 69634 5906 69646
rect 5854 69570 5906 69582
rect 6190 69634 6242 69646
rect 6190 69570 6242 69582
rect 6302 69634 6354 69646
rect 6302 69570 6354 69582
rect 28142 69634 28194 69646
rect 28142 69570 28194 69582
rect 31726 69634 31778 69646
rect 31726 69570 31778 69582
rect 32734 69634 32786 69646
rect 32734 69570 32786 69582
rect 33518 69634 33570 69646
rect 33518 69570 33570 69582
rect 1934 69522 1986 69534
rect 1934 69458 1986 69470
rect 3166 69522 3218 69534
rect 3166 69458 3218 69470
rect 4174 69522 4226 69534
rect 4174 69458 4226 69470
rect 4510 69522 4562 69534
rect 4510 69458 4562 69470
rect 4958 69522 5010 69534
rect 4958 69458 5010 69470
rect 7198 69522 7250 69534
rect 34526 69522 34578 69534
rect 13682 69470 13694 69522
rect 13746 69470 13758 69522
rect 17154 69470 17166 69522
rect 17218 69470 17230 69522
rect 19282 69470 19294 69522
rect 19346 69470 19358 69522
rect 22978 69470 22990 69522
rect 23042 69470 23054 69522
rect 25106 69470 25118 69522
rect 25170 69470 25182 69522
rect 7198 69458 7250 69470
rect 34526 69458 34578 69470
rect 34862 69522 34914 69534
rect 34862 69458 34914 69470
rect 35310 69522 35362 69534
rect 35310 69458 35362 69470
rect 35758 69522 35810 69534
rect 35758 69458 35810 69470
rect 3726 69410 3778 69422
rect 3726 69346 3778 69358
rect 5966 69410 6018 69422
rect 5966 69346 6018 69358
rect 7646 69410 7698 69422
rect 7646 69346 7698 69358
rect 7870 69410 7922 69422
rect 12462 69410 12514 69422
rect 8194 69358 8206 69410
rect 8258 69358 8270 69410
rect 9538 69358 9550 69410
rect 9602 69358 9614 69410
rect 10322 69358 10334 69410
rect 10386 69358 10398 69410
rect 7870 69346 7922 69358
rect 12462 69346 12514 69358
rect 13022 69410 13074 69422
rect 26126 69410 26178 69422
rect 27134 69410 27186 69422
rect 16594 69358 16606 69410
rect 16658 69358 16670 69410
rect 19954 69358 19966 69410
rect 20018 69358 20030 69410
rect 22194 69358 22206 69410
rect 22258 69358 22270 69410
rect 26786 69358 26798 69410
rect 26850 69358 26862 69410
rect 13022 69346 13074 69358
rect 26126 69346 26178 69358
rect 27134 69346 27186 69358
rect 28030 69410 28082 69422
rect 28030 69346 28082 69358
rect 28366 69410 28418 69422
rect 28366 69346 28418 69358
rect 28590 69410 28642 69422
rect 30158 69410 30210 69422
rect 33406 69410 33458 69422
rect 28802 69358 28814 69410
rect 28866 69358 28878 69410
rect 32050 69358 32062 69410
rect 32114 69358 32126 69410
rect 28590 69346 28642 69358
rect 30158 69346 30210 69358
rect 33406 69346 33458 69358
rect 34078 69410 34130 69422
rect 34078 69346 34130 69358
rect 11566 69298 11618 69310
rect 9090 69246 9102 69298
rect 9154 69246 9166 69298
rect 11566 69234 11618 69246
rect 11678 69298 11730 69310
rect 20526 69298 20578 69310
rect 15810 69246 15822 69298
rect 15874 69246 15886 69298
rect 11678 69234 11730 69246
rect 20526 69234 20578 69246
rect 20750 69298 20802 69310
rect 30046 69298 30098 69310
rect 20750 69234 20802 69246
rect 20862 69242 20914 69254
rect 2382 69186 2434 69198
rect 2382 69122 2434 69134
rect 2830 69186 2882 69198
rect 11902 69186 11954 69198
rect 10882 69134 10894 69186
rect 10946 69134 10958 69186
rect 2830 69122 2882 69134
rect 11902 69122 11954 69134
rect 12350 69186 12402 69198
rect 12350 69122 12402 69134
rect 12574 69186 12626 69198
rect 30046 69234 30098 69246
rect 30830 69298 30882 69310
rect 30830 69234 30882 69246
rect 32846 69242 32898 69254
rect 20862 69178 20914 69190
rect 21758 69186 21810 69198
rect 12574 69122 12626 69134
rect 21758 69122 21810 69134
rect 25790 69186 25842 69198
rect 25790 69122 25842 69134
rect 26014 69186 26066 69198
rect 26014 69122 26066 69134
rect 26238 69186 26290 69198
rect 26238 69122 26290 69134
rect 27246 69186 27298 69198
rect 27246 69122 27298 69134
rect 27358 69186 27410 69198
rect 27358 69122 27410 69134
rect 29710 69186 29762 69198
rect 29710 69122 29762 69134
rect 29934 69186 29986 69198
rect 29934 69122 29986 69134
rect 30718 69186 30770 69198
rect 30718 69122 30770 69134
rect 31838 69186 31890 69198
rect 31838 69122 31890 69134
rect 32734 69186 32786 69198
rect 32846 69178 32898 69190
rect 36206 69186 36258 69198
rect 32734 69122 32786 69134
rect 36206 69122 36258 69134
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 5070 68850 5122 68862
rect 5070 68786 5122 68798
rect 9886 68850 9938 68862
rect 9886 68786 9938 68798
rect 18510 68850 18562 68862
rect 18510 68786 18562 68798
rect 24894 68850 24946 68862
rect 24894 68786 24946 68798
rect 26014 68850 26066 68862
rect 26014 68786 26066 68798
rect 26126 68850 26178 68862
rect 26126 68786 26178 68798
rect 32958 68850 33010 68862
rect 32958 68786 33010 68798
rect 33966 68850 34018 68862
rect 33966 68786 34018 68798
rect 4398 68738 4450 68750
rect 4398 68674 4450 68686
rect 9774 68738 9826 68750
rect 25678 68738 25730 68750
rect 32846 68738 32898 68750
rect 21186 68686 21198 68738
rect 21250 68686 21262 68738
rect 30034 68686 30046 68738
rect 30098 68686 30110 68738
rect 9774 68674 9826 68686
rect 25678 68674 25730 68686
rect 32846 68674 32898 68686
rect 33518 68738 33570 68750
rect 33518 68674 33570 68686
rect 2046 68626 2098 68638
rect 2046 68562 2098 68574
rect 2382 68626 2434 68638
rect 18174 68626 18226 68638
rect 8866 68574 8878 68626
rect 8930 68574 8942 68626
rect 10434 68574 10446 68626
rect 10498 68574 10510 68626
rect 16706 68574 16718 68626
rect 16770 68574 16782 68626
rect 2382 68562 2434 68574
rect 18174 68562 18226 68574
rect 18398 68626 18450 68638
rect 25902 68626 25954 68638
rect 19170 68574 19182 68626
rect 19234 68574 19246 68626
rect 18398 68562 18450 68574
rect 25902 68562 25954 68574
rect 26238 68626 26290 68638
rect 26238 68562 26290 68574
rect 27246 68626 27298 68638
rect 27246 68562 27298 68574
rect 27470 68626 27522 68638
rect 27470 68562 27522 68574
rect 28254 68626 28306 68638
rect 28254 68562 28306 68574
rect 29038 68626 29090 68638
rect 32286 68626 32338 68638
rect 31602 68574 31614 68626
rect 31666 68574 31678 68626
rect 32610 68574 32622 68626
rect 32674 68574 32686 68626
rect 29038 68562 29090 68574
rect 32286 68562 32338 68574
rect 2942 68514 2994 68526
rect 2942 68450 2994 68462
rect 3390 68514 3442 68526
rect 3390 68450 3442 68462
rect 3838 68514 3890 68526
rect 3838 68450 3890 68462
rect 5182 68514 5234 68526
rect 5182 68450 5234 68462
rect 6078 68514 6130 68526
rect 28702 68514 28754 68526
rect 34414 68514 34466 68526
rect 8194 68462 8206 68514
rect 8258 68462 8270 68514
rect 11778 68462 11790 68514
rect 11842 68462 11854 68514
rect 31378 68462 31390 68514
rect 31442 68462 31454 68514
rect 6078 68450 6130 68462
rect 28702 68450 28754 68462
rect 34414 68450 34466 68462
rect 34862 68514 34914 68526
rect 34862 68450 34914 68462
rect 35310 68514 35362 68526
rect 35310 68450 35362 68462
rect 4286 68402 4338 68414
rect 4286 68338 4338 68350
rect 5294 68402 5346 68414
rect 5294 68338 5346 68350
rect 10670 68402 10722 68414
rect 10670 68338 10722 68350
rect 10894 68402 10946 68414
rect 10894 68338 10946 68350
rect 11006 68402 11058 68414
rect 11006 68338 11058 68350
rect 18510 68402 18562 68414
rect 26898 68350 26910 68402
rect 26962 68350 26974 68402
rect 29922 68350 29934 68402
rect 29986 68350 29998 68402
rect 30930 68350 30942 68402
rect 30994 68350 31006 68402
rect 18510 68338 18562 68350
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 12462 68066 12514 68078
rect 5506 68014 5518 68066
rect 5570 68063 5582 68066
rect 5730 68063 5742 68066
rect 5570 68017 5742 68063
rect 5570 68014 5582 68017
rect 5730 68014 5742 68017
rect 5794 68014 5806 68066
rect 12462 68002 12514 68014
rect 12798 68066 12850 68078
rect 12798 68002 12850 68014
rect 12910 68066 12962 68078
rect 12910 68002 12962 68014
rect 14030 68066 14082 68078
rect 14030 68002 14082 68014
rect 29598 68066 29650 68078
rect 29598 68002 29650 68014
rect 31726 68066 31778 68078
rect 31726 68002 31778 68014
rect 3726 67954 3778 67966
rect 3726 67890 3778 67902
rect 7198 67954 7250 67966
rect 7198 67890 7250 67902
rect 7982 67954 8034 67966
rect 7982 67890 8034 67902
rect 10222 67954 10274 67966
rect 10222 67890 10274 67902
rect 11678 67954 11730 67966
rect 11678 67890 11730 67902
rect 13806 67954 13858 67966
rect 17166 67954 17218 67966
rect 23550 67954 23602 67966
rect 28814 67954 28866 67966
rect 15698 67902 15710 67954
rect 15762 67902 15774 67954
rect 17826 67902 17838 67954
rect 17890 67902 17902 67954
rect 20066 67902 20078 67954
rect 20130 67902 20142 67954
rect 26002 67902 26014 67954
rect 26066 67902 26078 67954
rect 28130 67902 28142 67954
rect 28194 67902 28206 67954
rect 13806 67890 13858 67902
rect 17166 67890 17218 67902
rect 23550 67890 23602 67902
rect 28814 67890 28866 67902
rect 2830 67842 2882 67854
rect 2830 67778 2882 67790
rect 4174 67842 4226 67854
rect 4174 67778 4226 67790
rect 4622 67842 4674 67854
rect 4622 67778 4674 67790
rect 5966 67842 6018 67854
rect 5966 67778 6018 67790
rect 8430 67842 8482 67854
rect 8430 67778 8482 67790
rect 9326 67842 9378 67854
rect 9326 67778 9378 67790
rect 10110 67842 10162 67854
rect 10110 67778 10162 67790
rect 10334 67842 10386 67854
rect 10334 67778 10386 67790
rect 11454 67842 11506 67854
rect 11454 67778 11506 67790
rect 12574 67842 12626 67854
rect 12574 67778 12626 67790
rect 14254 67842 14306 67854
rect 21758 67842 21810 67854
rect 23438 67842 23490 67854
rect 14466 67790 14478 67842
rect 14530 67790 14542 67842
rect 15586 67790 15598 67842
rect 15650 67790 15662 67842
rect 16258 67790 16270 67842
rect 16322 67790 16334 67842
rect 20738 67790 20750 67842
rect 20802 67790 20814 67842
rect 22082 67790 22094 67842
rect 22146 67790 22158 67842
rect 14254 67778 14306 67790
rect 21758 67778 21810 67790
rect 23438 67778 23490 67790
rect 23662 67842 23714 67854
rect 24446 67842 24498 67854
rect 23874 67790 23886 67842
rect 23938 67790 23950 67842
rect 23662 67778 23714 67790
rect 24446 67778 24498 67790
rect 24782 67842 24834 67854
rect 30718 67842 30770 67854
rect 25330 67790 25342 67842
rect 25394 67790 25406 67842
rect 24782 67778 24834 67790
rect 30718 67778 30770 67790
rect 31614 67842 31666 67854
rect 31614 67778 31666 67790
rect 32398 67842 32450 67854
rect 32398 67778 32450 67790
rect 32734 67842 32786 67854
rect 32734 67778 32786 67790
rect 3278 67730 3330 67742
rect 3278 67666 3330 67678
rect 7870 67730 7922 67742
rect 7870 67666 7922 67678
rect 8206 67730 8258 67742
rect 8206 67666 8258 67678
rect 8990 67730 9042 67742
rect 8990 67666 9042 67678
rect 9550 67730 9602 67742
rect 9550 67666 9602 67678
rect 10558 67730 10610 67742
rect 10558 67666 10610 67678
rect 11230 67730 11282 67742
rect 11230 67666 11282 67678
rect 11790 67730 11842 67742
rect 21646 67730 21698 67742
rect 15698 67678 15710 67730
rect 15762 67678 15774 67730
rect 16594 67678 16606 67730
rect 16658 67678 16670 67730
rect 11790 67666 11842 67678
rect 21646 67666 21698 67678
rect 23214 67730 23266 67742
rect 23214 67666 23266 67678
rect 29934 67730 29986 67742
rect 29934 67666 29986 67678
rect 30606 67730 30658 67742
rect 30606 67666 30658 67678
rect 31726 67730 31778 67742
rect 31726 67666 31778 67678
rect 33966 67730 34018 67742
rect 33966 67666 34018 67678
rect 1934 67618 1986 67630
rect 1934 67554 1986 67566
rect 2382 67618 2434 67630
rect 2382 67554 2434 67566
rect 4958 67618 5010 67630
rect 4958 67554 5010 67566
rect 6078 67618 6130 67630
rect 6078 67554 6130 67566
rect 6302 67618 6354 67630
rect 6302 67554 6354 67566
rect 6862 67618 6914 67630
rect 6862 67554 6914 67566
rect 7086 67618 7138 67630
rect 7086 67554 7138 67566
rect 7310 67618 7362 67630
rect 7310 67554 7362 67566
rect 9102 67618 9154 67630
rect 9102 67554 9154 67566
rect 14366 67618 14418 67630
rect 14366 67554 14418 67566
rect 24558 67618 24610 67630
rect 24558 67554 24610 67566
rect 29710 67618 29762 67630
rect 29710 67554 29762 67566
rect 30382 67618 30434 67630
rect 30382 67554 30434 67566
rect 32510 67618 32562 67630
rect 32510 67554 32562 67566
rect 33070 67618 33122 67630
rect 33070 67554 33122 67566
rect 33518 67618 33570 67630
rect 33518 67554 33570 67566
rect 34414 67618 34466 67630
rect 34414 67554 34466 67566
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 3614 67282 3666 67294
rect 3614 67218 3666 67230
rect 6638 67282 6690 67294
rect 6638 67218 6690 67230
rect 8878 67282 8930 67294
rect 8878 67218 8930 67230
rect 17950 67282 18002 67294
rect 17950 67218 18002 67230
rect 31390 67282 31442 67294
rect 31390 67218 31442 67230
rect 31614 67282 31666 67294
rect 31614 67218 31666 67230
rect 31950 67282 32002 67294
rect 31950 67218 32002 67230
rect 3166 67170 3218 67182
rect 5406 67170 5458 67182
rect 4834 67118 4846 67170
rect 4898 67118 4910 67170
rect 3166 67106 3218 67118
rect 4622 67058 4674 67070
rect 4622 66994 4674 67006
rect 1934 66946 1986 66958
rect 1934 66882 1986 66894
rect 2382 66946 2434 66958
rect 2382 66882 2434 66894
rect 2718 66946 2770 66958
rect 2718 66882 2770 66894
rect 4174 66946 4226 66958
rect 4174 66882 4226 66894
rect 3378 66782 3390 66834
rect 3442 66831 3454 66834
rect 4849 66831 4895 67118
rect 5406 67106 5458 67118
rect 7422 67170 7474 67182
rect 7422 67106 7474 67118
rect 10110 67170 10162 67182
rect 10110 67106 10162 67118
rect 14926 67170 14978 67182
rect 22654 67170 22706 67182
rect 20066 67118 20078 67170
rect 20130 67118 20142 67170
rect 14926 67106 14978 67118
rect 22654 67106 22706 67118
rect 24334 67170 24386 67182
rect 24334 67106 24386 67118
rect 26126 67170 26178 67182
rect 26126 67106 26178 67118
rect 26238 67170 26290 67182
rect 26238 67106 26290 67118
rect 26910 67170 26962 67182
rect 26910 67106 26962 67118
rect 27134 67170 27186 67182
rect 27134 67106 27186 67118
rect 28590 67170 28642 67182
rect 32398 67170 32450 67182
rect 29362 67118 29374 67170
rect 29426 67118 29438 67170
rect 28590 67106 28642 67118
rect 32398 67106 32450 67118
rect 32846 67170 32898 67182
rect 32846 67106 32898 67118
rect 10334 67058 10386 67070
rect 6962 67006 6974 67058
rect 7026 67055 7038 67058
rect 7186 67055 7198 67058
rect 7026 67009 7198 67055
rect 7026 67006 7038 67009
rect 7186 67006 7198 67009
rect 7250 67006 7262 67058
rect 7634 67006 7646 67058
rect 7698 67006 7710 67058
rect 8754 67006 8766 67058
rect 8818 67006 8830 67058
rect 10334 66994 10386 67006
rect 10558 67058 10610 67070
rect 15150 67058 15202 67070
rect 11554 67006 11566 67058
rect 11618 67006 11630 67058
rect 10558 66994 10610 67006
rect 15150 66994 15202 67006
rect 15598 67058 15650 67070
rect 18286 67058 18338 67070
rect 26014 67058 26066 67070
rect 16594 67006 16606 67058
rect 16658 67006 16670 67058
rect 18498 67006 18510 67058
rect 18562 67006 18574 67058
rect 19282 67006 19294 67058
rect 19346 67006 19358 67058
rect 23874 67006 23886 67058
rect 23938 67006 23950 67058
rect 25666 67006 25678 67058
rect 25730 67006 25742 67058
rect 15598 66994 15650 67006
rect 18286 66994 18338 67006
rect 26014 66994 26066 67006
rect 26798 67058 26850 67070
rect 31278 67058 31330 67070
rect 27906 67006 27918 67058
rect 27970 67006 27982 67058
rect 29586 67006 29598 67058
rect 29650 67006 29662 67058
rect 30258 67006 30270 67058
rect 30322 67006 30334 67058
rect 30594 67006 30606 67058
rect 30658 67006 30670 67058
rect 26798 66994 26850 67006
rect 31278 66994 31330 67006
rect 4958 66946 5010 66958
rect 4958 66882 5010 66894
rect 5854 66946 5906 66958
rect 10446 66946 10498 66958
rect 15374 66946 15426 66958
rect 6626 66894 6638 66946
rect 6690 66894 6702 66946
rect 8530 66894 8542 66946
rect 8594 66894 8606 66946
rect 12226 66894 12238 66946
rect 12290 66894 12302 66946
rect 14354 66894 14366 66946
rect 14418 66894 14430 66946
rect 5854 66882 5906 66894
rect 10446 66882 10498 66894
rect 15374 66882 15426 66894
rect 16942 66946 16994 66958
rect 16942 66882 16994 66894
rect 17838 66946 17890 66958
rect 24894 66946 24946 66958
rect 22194 66894 22206 66946
rect 22258 66894 22270 66946
rect 23986 66894 23998 66946
rect 24050 66894 24062 66946
rect 27794 66894 27806 66946
rect 27858 66894 27870 66946
rect 29250 66894 29262 66946
rect 29314 66894 29326 66946
rect 17838 66882 17890 66894
rect 24894 66882 24946 66894
rect 3442 66785 4895 66831
rect 6414 66834 6466 66846
rect 3442 66782 3454 66785
rect 6414 66770 6466 66782
rect 7310 66834 7362 66846
rect 7310 66770 7362 66782
rect 16046 66834 16098 66846
rect 16046 66770 16098 66782
rect 16606 66834 16658 66846
rect 16606 66770 16658 66782
rect 18062 66834 18114 66846
rect 18062 66770 18114 66782
rect 27582 66834 27634 66846
rect 32050 66782 32062 66834
rect 32114 66831 32126 66834
rect 32610 66831 32622 66834
rect 32114 66785 32622 66831
rect 32114 66782 32126 66785
rect 32610 66782 32622 66785
rect 32674 66782 32686 66834
rect 27582 66770 27634 66782
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 8094 66498 8146 66510
rect 5954 66446 5966 66498
rect 6018 66495 6030 66498
rect 6402 66495 6414 66498
rect 6018 66449 6414 66495
rect 6018 66446 6030 66449
rect 6402 66446 6414 66449
rect 6466 66446 6478 66498
rect 8094 66434 8146 66446
rect 9326 66498 9378 66510
rect 29934 66498 29986 66510
rect 28802 66446 28814 66498
rect 28866 66446 28878 66498
rect 9326 66434 9378 66446
rect 29934 66434 29986 66446
rect 2158 66386 2210 66398
rect 2158 66322 2210 66334
rect 2606 66386 2658 66398
rect 2606 66322 2658 66334
rect 4062 66386 4114 66398
rect 4062 66322 4114 66334
rect 4622 66386 4674 66398
rect 4622 66322 4674 66334
rect 6302 66386 6354 66398
rect 6302 66322 6354 66334
rect 6750 66386 6802 66398
rect 6750 66322 6802 66334
rect 9214 66386 9266 66398
rect 9214 66322 9266 66334
rect 11902 66386 11954 66398
rect 19294 66386 19346 66398
rect 20862 66386 20914 66398
rect 13682 66334 13694 66386
rect 13746 66334 13758 66386
rect 20066 66334 20078 66386
rect 20130 66334 20142 66386
rect 11902 66322 11954 66334
rect 19294 66322 19346 66334
rect 20862 66322 20914 66334
rect 22878 66386 22930 66398
rect 30606 66386 30658 66398
rect 32062 66386 32114 66398
rect 23426 66334 23438 66386
rect 23490 66334 23502 66386
rect 29586 66334 29598 66386
rect 29650 66334 29662 66386
rect 31490 66334 31502 66386
rect 31554 66334 31566 66386
rect 22878 66322 22930 66334
rect 30606 66322 30658 66334
rect 32062 66322 32114 66334
rect 12686 66274 12738 66286
rect 18510 66274 18562 66286
rect 22766 66274 22818 66286
rect 26910 66274 26962 66286
rect 3154 66222 3166 66274
rect 3218 66222 3230 66274
rect 10546 66222 10558 66274
rect 10610 66222 10622 66274
rect 16482 66222 16494 66274
rect 16546 66222 16558 66274
rect 17154 66222 17166 66274
rect 17218 66222 17230 66274
rect 19954 66222 19966 66274
rect 20018 66222 20030 66274
rect 22194 66222 22206 66274
rect 22258 66222 22270 66274
rect 26226 66222 26238 66274
rect 26290 66222 26302 66274
rect 12686 66210 12738 66222
rect 18510 66210 18562 66222
rect 22766 66210 22818 66222
rect 26910 66210 26962 66222
rect 27134 66274 27186 66286
rect 27134 66210 27186 66222
rect 27582 66274 27634 66286
rect 27582 66210 27634 66222
rect 28254 66274 28306 66286
rect 31266 66222 31278 66274
rect 31330 66222 31342 66274
rect 28254 66210 28306 66222
rect 3390 66162 3442 66174
rect 3390 66098 3442 66110
rect 6862 66162 6914 66174
rect 6862 66098 6914 66110
rect 7422 66162 7474 66174
rect 7422 66098 7474 66110
rect 8318 66162 8370 66174
rect 17390 66162 17442 66174
rect 11554 66110 11566 66162
rect 11618 66110 11630 66162
rect 15810 66110 15822 66162
rect 15874 66110 15886 66162
rect 8318 66098 8370 66110
rect 17390 66098 17442 66110
rect 17502 66162 17554 66174
rect 17502 66098 17554 66110
rect 18622 66162 18674 66174
rect 28142 66162 28194 66174
rect 25554 66110 25566 66162
rect 25618 66110 25630 66162
rect 18622 66098 18674 66110
rect 28142 66098 28194 66110
rect 28366 66162 28418 66174
rect 28366 66098 28418 66110
rect 29710 66162 29762 66174
rect 29710 66098 29762 66110
rect 5070 66050 5122 66062
rect 5070 65986 5122 65998
rect 5742 66050 5794 66062
rect 5742 65986 5794 65998
rect 7534 66050 7586 66062
rect 7534 65986 7586 65998
rect 8206 66050 8258 66062
rect 8206 65986 8258 65998
rect 9102 66050 9154 66062
rect 12798 66050 12850 66062
rect 9986 65998 9998 66050
rect 10050 65998 10062 66050
rect 9102 65986 9154 65998
rect 12798 65986 12850 65998
rect 13022 66050 13074 66062
rect 18846 66050 18898 66062
rect 17938 65998 17950 66050
rect 18002 65998 18014 66050
rect 13022 65986 13074 65998
rect 18846 65986 18898 65998
rect 27022 66050 27074 66062
rect 27022 65986 27074 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 8094 65714 8146 65726
rect 7422 65658 7474 65670
rect 4846 65602 4898 65614
rect 8094 65650 8146 65662
rect 8318 65714 8370 65726
rect 8318 65650 8370 65662
rect 16382 65714 16434 65726
rect 16382 65650 16434 65662
rect 18174 65714 18226 65726
rect 18174 65650 18226 65662
rect 21534 65714 21586 65726
rect 21534 65650 21586 65662
rect 21646 65714 21698 65726
rect 21646 65650 21698 65662
rect 21758 65714 21810 65726
rect 21758 65650 21810 65662
rect 21870 65714 21922 65726
rect 21870 65650 21922 65662
rect 24894 65714 24946 65726
rect 24894 65650 24946 65662
rect 30494 65714 30546 65726
rect 30494 65650 30546 65662
rect 31054 65714 31106 65726
rect 31054 65650 31106 65662
rect 7422 65594 7474 65606
rect 8206 65602 8258 65614
rect 4846 65538 4898 65550
rect 7310 65546 7362 65558
rect 2270 65490 2322 65502
rect 2270 65426 2322 65438
rect 4062 65490 4114 65502
rect 4062 65426 4114 65438
rect 5406 65490 5458 65502
rect 8206 65538 8258 65550
rect 10222 65602 10274 65614
rect 16270 65602 16322 65614
rect 12450 65550 12462 65602
rect 12514 65550 12526 65602
rect 10222 65538 10274 65550
rect 16270 65538 16322 65550
rect 17726 65602 17778 65614
rect 17726 65538 17778 65550
rect 18622 65602 18674 65614
rect 18622 65538 18674 65550
rect 20190 65602 20242 65614
rect 20190 65538 20242 65550
rect 20302 65602 20354 65614
rect 20302 65538 20354 65550
rect 21310 65602 21362 65614
rect 21310 65538 21362 65550
rect 22542 65602 22594 65614
rect 26686 65602 26738 65614
rect 30606 65602 30658 65614
rect 23538 65550 23550 65602
rect 23602 65550 23614 65602
rect 23874 65550 23886 65602
rect 23938 65550 23950 65602
rect 27346 65550 27358 65602
rect 27410 65550 27422 65602
rect 27906 65550 27918 65602
rect 27970 65550 27982 65602
rect 22542 65538 22594 65550
rect 26686 65538 26738 65550
rect 30606 65538 30658 65550
rect 7310 65482 7362 65494
rect 7646 65490 7698 65502
rect 5406 65426 5458 65438
rect 7646 65426 7698 65438
rect 8766 65490 8818 65502
rect 15598 65490 15650 65502
rect 11218 65438 11230 65490
rect 11282 65438 11294 65490
rect 13794 65438 13806 65490
rect 13858 65438 13870 65490
rect 14802 65438 14814 65490
rect 14866 65438 14878 65490
rect 8766 65426 8818 65438
rect 15598 65426 15650 65438
rect 16606 65490 16658 65502
rect 16606 65426 16658 65438
rect 16718 65490 16770 65502
rect 16718 65426 16770 65438
rect 17950 65490 18002 65502
rect 17950 65426 18002 65438
rect 18286 65490 18338 65502
rect 18286 65426 18338 65438
rect 19182 65490 19234 65502
rect 23438 65490 23490 65502
rect 22754 65438 22766 65490
rect 22818 65438 22830 65490
rect 19182 65426 19234 65438
rect 23438 65426 23490 65438
rect 24222 65490 24274 65502
rect 29710 65490 29762 65502
rect 26002 65438 26014 65490
rect 26066 65438 26078 65490
rect 26450 65438 26462 65490
rect 26514 65438 26526 65490
rect 27682 65438 27694 65490
rect 27746 65438 27758 65490
rect 29474 65438 29486 65490
rect 29538 65438 29550 65490
rect 24222 65426 24274 65438
rect 29710 65426 29762 65438
rect 30270 65490 30322 65502
rect 30270 65426 30322 65438
rect 1822 65378 1874 65390
rect 1822 65314 1874 65326
rect 2718 65378 2770 65390
rect 2718 65314 2770 65326
rect 3054 65378 3106 65390
rect 3054 65314 3106 65326
rect 3614 65378 3666 65390
rect 3614 65314 3666 65326
rect 4510 65378 4562 65390
rect 4510 65314 4562 65326
rect 6302 65378 6354 65390
rect 6302 65314 6354 65326
rect 6750 65378 6802 65390
rect 28814 65378 28866 65390
rect 11106 65326 11118 65378
rect 11170 65326 11182 65378
rect 13458 65326 13470 65378
rect 13522 65326 13534 65378
rect 16258 65326 16270 65378
rect 16322 65326 16334 65378
rect 6750 65314 6802 65326
rect 28814 65314 28866 65326
rect 5518 65266 5570 65278
rect 10110 65266 10162 65278
rect 4498 65214 4510 65266
rect 4562 65263 4574 65266
rect 5170 65263 5182 65266
rect 4562 65217 5182 65263
rect 4562 65214 4574 65217
rect 5170 65214 5182 65217
rect 5234 65214 5246 65266
rect 6514 65214 6526 65266
rect 6578 65263 6590 65266
rect 7074 65263 7086 65266
rect 6578 65217 7086 65263
rect 6578 65214 6590 65217
rect 7074 65214 7086 65217
rect 7138 65214 7150 65266
rect 5518 65202 5570 65214
rect 10110 65202 10162 65214
rect 10446 65266 10498 65278
rect 10446 65202 10498 65214
rect 18174 65266 18226 65278
rect 18174 65202 18226 65214
rect 19742 65266 19794 65278
rect 19742 65202 19794 65214
rect 19966 65266 20018 65278
rect 19966 65202 20018 65214
rect 20526 65266 20578 65278
rect 20526 65202 20578 65214
rect 24446 65266 24498 65278
rect 24446 65202 24498 65214
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 11902 64930 11954 64942
rect 15374 64930 15426 64942
rect 2034 64878 2046 64930
rect 2098 64927 2110 64930
rect 2594 64927 2606 64930
rect 2098 64881 2606 64927
rect 2098 64878 2110 64881
rect 2594 64878 2606 64881
rect 2658 64878 2670 64930
rect 3602 64878 3614 64930
rect 3666 64927 3678 64930
rect 3666 64881 4895 64927
rect 3666 64878 3678 64881
rect 1934 64818 1986 64830
rect 1934 64754 1986 64766
rect 2382 64818 2434 64830
rect 2382 64754 2434 64766
rect 3166 64706 3218 64718
rect 3166 64642 3218 64654
rect 3614 64706 3666 64718
rect 4849 64706 4895 64881
rect 14242 64878 14254 64930
rect 14306 64878 14318 64930
rect 11902 64866 11954 64878
rect 15374 64866 15426 64878
rect 16046 64930 16098 64942
rect 16046 64866 16098 64878
rect 27022 64930 27074 64942
rect 27022 64866 27074 64878
rect 4958 64818 5010 64830
rect 17726 64818 17778 64830
rect 22094 64818 22146 64830
rect 6066 64766 6078 64818
rect 6130 64766 6142 64818
rect 14018 64766 14030 64818
rect 14082 64766 14094 64818
rect 20514 64766 20526 64818
rect 20578 64766 20590 64818
rect 4958 64754 5010 64766
rect 17726 64754 17778 64766
rect 22094 64754 22146 64766
rect 23102 64818 23154 64830
rect 23102 64754 23154 64766
rect 23998 64818 24050 64830
rect 23998 64754 24050 64766
rect 27470 64818 27522 64830
rect 29822 64818 29874 64830
rect 28242 64766 28254 64818
rect 28306 64766 28318 64818
rect 27470 64754 27522 64766
rect 29822 64754 29874 64766
rect 30270 64818 30322 64830
rect 30270 64754 30322 64766
rect 9438 64706 9490 64718
rect 15486 64706 15538 64718
rect 4834 64654 4846 64706
rect 4898 64654 4910 64706
rect 7522 64654 7534 64706
rect 7586 64654 7598 64706
rect 14354 64654 14366 64706
rect 14418 64654 14430 64706
rect 3614 64642 3666 64654
rect 9438 64642 9490 64654
rect 15486 64642 15538 64654
rect 15710 64706 15762 64718
rect 15710 64642 15762 64654
rect 15934 64706 15986 64718
rect 15934 64642 15986 64654
rect 16830 64706 16882 64718
rect 18958 64706 19010 64718
rect 23774 64706 23826 64718
rect 17154 64654 17166 64706
rect 17218 64654 17230 64706
rect 19842 64654 19854 64706
rect 19906 64654 19918 64706
rect 20178 64654 20190 64706
rect 20242 64654 20254 64706
rect 16830 64642 16882 64654
rect 18958 64642 19010 64654
rect 23774 64642 23826 64654
rect 23886 64706 23938 64718
rect 23886 64642 23938 64654
rect 24110 64706 24162 64718
rect 25118 64706 25170 64718
rect 24322 64654 24334 64706
rect 24386 64654 24398 64706
rect 24110 64642 24162 64654
rect 25118 64642 25170 64654
rect 25342 64706 25394 64718
rect 25342 64642 25394 64654
rect 26350 64706 26402 64718
rect 26674 64654 26686 64706
rect 26738 64654 26750 64706
rect 28018 64654 28030 64706
rect 28082 64654 28094 64706
rect 26350 64642 26402 64654
rect 2830 64594 2882 64606
rect 2830 64530 2882 64542
rect 4510 64594 4562 64606
rect 9662 64594 9714 64606
rect 6514 64542 6526 64594
rect 6578 64542 6590 64594
rect 4510 64530 4562 64542
rect 9662 64530 9714 64542
rect 9774 64594 9826 64606
rect 18398 64594 18450 64606
rect 9986 64542 9998 64594
rect 10050 64542 10062 64594
rect 12114 64542 12126 64594
rect 12178 64542 12190 64594
rect 12562 64542 12574 64594
rect 12626 64542 12638 64594
rect 9774 64530 9826 64542
rect 18398 64530 18450 64542
rect 25678 64594 25730 64606
rect 25678 64530 25730 64542
rect 26910 64594 26962 64606
rect 26910 64530 26962 64542
rect 4062 64482 4114 64494
rect 8990 64482 9042 64494
rect 7858 64430 7870 64482
rect 7922 64430 7934 64482
rect 4062 64418 4114 64430
rect 8990 64418 9042 64430
rect 9550 64482 9602 64494
rect 9550 64418 9602 64430
rect 10894 64482 10946 64494
rect 10894 64418 10946 64430
rect 11566 64482 11618 64494
rect 11566 64418 11618 64430
rect 18286 64482 18338 64494
rect 18286 64418 18338 64430
rect 18510 64482 18562 64494
rect 18510 64418 18562 64430
rect 20862 64482 20914 64494
rect 20862 64418 20914 64430
rect 21982 64482 22034 64494
rect 21982 64418 22034 64430
rect 22206 64482 22258 64494
rect 22206 64418 22258 64430
rect 22430 64482 22482 64494
rect 22430 64418 22482 64430
rect 25566 64482 25618 64494
rect 25566 64418 25618 64430
rect 25790 64482 25842 64494
rect 25790 64418 25842 64430
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 1934 64146 1986 64158
rect 1934 64082 1986 64094
rect 2718 64146 2770 64158
rect 2718 64082 2770 64094
rect 4622 64146 4674 64158
rect 4622 64082 4674 64094
rect 5518 64146 5570 64158
rect 5518 64082 5570 64094
rect 5854 64146 5906 64158
rect 5854 64082 5906 64094
rect 7198 64146 7250 64158
rect 11454 64146 11506 64158
rect 8194 64094 8206 64146
rect 8258 64094 8270 64146
rect 7198 64082 7250 64094
rect 11454 64082 11506 64094
rect 12126 64146 12178 64158
rect 12126 64082 12178 64094
rect 15038 64146 15090 64158
rect 15038 64082 15090 64094
rect 15150 64146 15202 64158
rect 15150 64082 15202 64094
rect 15262 64146 15314 64158
rect 15262 64082 15314 64094
rect 16382 64146 16434 64158
rect 16382 64082 16434 64094
rect 16494 64146 16546 64158
rect 16494 64082 16546 64094
rect 16606 64146 16658 64158
rect 16606 64082 16658 64094
rect 18174 64146 18226 64158
rect 18174 64082 18226 64094
rect 19182 64146 19234 64158
rect 19182 64082 19234 64094
rect 20302 64146 20354 64158
rect 20302 64082 20354 64094
rect 20526 64146 20578 64158
rect 20526 64082 20578 64094
rect 22766 64146 22818 64158
rect 22766 64082 22818 64094
rect 24110 64146 24162 64158
rect 24110 64082 24162 64094
rect 24894 64146 24946 64158
rect 24894 64082 24946 64094
rect 26798 64146 26850 64158
rect 26798 64082 26850 64094
rect 27806 64146 27858 64158
rect 27806 64082 27858 64094
rect 28590 64146 28642 64158
rect 28590 64082 28642 64094
rect 28926 64146 28978 64158
rect 28926 64082 28978 64094
rect 12350 64034 12402 64046
rect 12350 63970 12402 63982
rect 19070 64034 19122 64046
rect 19070 63970 19122 63982
rect 19630 64034 19682 64046
rect 19630 63970 19682 63982
rect 20190 64034 20242 64046
rect 20190 63970 20242 63982
rect 23326 64034 23378 64046
rect 23326 63970 23378 63982
rect 25790 64034 25842 64046
rect 25790 63970 25842 63982
rect 25902 64034 25954 64046
rect 25902 63970 25954 63982
rect 2382 63922 2434 63934
rect 2382 63858 2434 63870
rect 3726 63922 3778 63934
rect 3726 63858 3778 63870
rect 6302 63922 6354 63934
rect 6302 63858 6354 63870
rect 6862 63922 6914 63934
rect 6862 63858 6914 63870
rect 8766 63922 8818 63934
rect 12014 63922 12066 63934
rect 9986 63870 9998 63922
rect 10050 63870 10062 63922
rect 8766 63858 8818 63870
rect 12014 63858 12066 63870
rect 12574 63922 12626 63934
rect 15486 63922 15538 63934
rect 18398 63922 18450 63934
rect 13570 63870 13582 63922
rect 13634 63870 13646 63922
rect 16930 63870 16942 63922
rect 16994 63870 17006 63922
rect 18050 63870 18062 63922
rect 18114 63870 18126 63922
rect 12574 63858 12626 63870
rect 15486 63858 15538 63870
rect 18398 63858 18450 63870
rect 19294 63922 19346 63934
rect 22206 63922 22258 63934
rect 21522 63870 21534 63922
rect 21586 63870 21598 63922
rect 19294 63858 19346 63870
rect 22206 63858 22258 63870
rect 25566 63922 25618 63934
rect 25566 63858 25618 63870
rect 26686 63922 26738 63934
rect 26686 63858 26738 63870
rect 26910 63922 26962 63934
rect 26910 63858 26962 63870
rect 27358 63922 27410 63934
rect 27358 63858 27410 63870
rect 3166 63810 3218 63822
rect 3166 63746 3218 63758
rect 4062 63810 4114 63822
rect 4062 63746 4114 63758
rect 4958 63810 5010 63822
rect 4958 63746 5010 63758
rect 7646 63810 7698 63822
rect 7646 63746 7698 63758
rect 10334 63810 10386 63822
rect 17726 63810 17778 63822
rect 13906 63758 13918 63810
rect 13970 63758 13982 63810
rect 10334 63746 10386 63758
rect 17726 63746 17778 63758
rect 18286 63810 18338 63822
rect 21298 63758 21310 63810
rect 21362 63758 21374 63810
rect 18286 63746 18338 63758
rect 8542 63698 8594 63710
rect 15710 63698 15762 63710
rect 1698 63646 1710 63698
rect 1762 63695 1774 63698
rect 2818 63695 2830 63698
rect 1762 63649 2830 63695
rect 1762 63646 1774 63649
rect 2818 63646 2830 63649
rect 2882 63646 2894 63698
rect 4050 63646 4062 63698
rect 4114 63695 4126 63698
rect 6850 63695 6862 63698
rect 4114 63649 6862 63695
rect 4114 63646 4126 63649
rect 6850 63646 6862 63649
rect 6914 63646 6926 63698
rect 13682 63646 13694 63698
rect 13746 63646 13758 63698
rect 8542 63634 8594 63646
rect 15710 63634 15762 63646
rect 23886 63698 23938 63710
rect 23886 63634 23938 63646
rect 24222 63698 24274 63710
rect 24222 63634 24274 63646
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 10334 63362 10386 63374
rect 19742 63362 19794 63374
rect 2482 63310 2494 63362
rect 2546 63359 2558 63362
rect 3266 63359 3278 63362
rect 2546 63313 3278 63359
rect 2546 63310 2558 63313
rect 3266 63310 3278 63313
rect 3330 63359 3342 63362
rect 4498 63359 4510 63362
rect 3330 63313 4510 63359
rect 3330 63310 3342 63313
rect 4498 63310 4510 63313
rect 4562 63310 4574 63362
rect 6514 63310 6526 63362
rect 6578 63359 6590 63362
rect 8642 63359 8654 63362
rect 6578 63313 8654 63359
rect 6578 63310 6590 63313
rect 8642 63310 8654 63313
rect 8706 63310 8718 63362
rect 15922 63310 15934 63362
rect 15986 63310 15998 63362
rect 10334 63298 10386 63310
rect 19742 63298 19794 63310
rect 22878 63362 22930 63374
rect 22878 63298 22930 63310
rect 24334 63362 24386 63374
rect 24334 63298 24386 63310
rect 25118 63362 25170 63374
rect 25118 63298 25170 63310
rect 1934 63250 1986 63262
rect 1934 63186 1986 63198
rect 2718 63250 2770 63262
rect 2718 63186 2770 63198
rect 3166 63250 3218 63262
rect 3166 63186 3218 63198
rect 3614 63250 3666 63262
rect 3614 63186 3666 63198
rect 4174 63250 4226 63262
rect 4174 63186 4226 63198
rect 4622 63250 4674 63262
rect 4622 63186 4674 63198
rect 6526 63250 6578 63262
rect 6526 63186 6578 63198
rect 6862 63250 6914 63262
rect 6862 63186 6914 63198
rect 8206 63250 8258 63262
rect 8206 63186 8258 63198
rect 9998 63250 10050 63262
rect 9998 63186 10050 63198
rect 10558 63250 10610 63262
rect 12910 63250 12962 63262
rect 12002 63198 12014 63250
rect 12066 63198 12078 63250
rect 10558 63186 10610 63198
rect 12910 63186 12962 63198
rect 15262 63250 15314 63262
rect 20414 63250 20466 63262
rect 16034 63198 16046 63250
rect 16098 63198 16110 63250
rect 17602 63198 17614 63250
rect 17666 63198 17678 63250
rect 18386 63198 18398 63250
rect 18450 63198 18462 63250
rect 15262 63186 15314 63198
rect 20414 63186 20466 63198
rect 22990 63250 23042 63262
rect 22990 63186 23042 63198
rect 23662 63250 23714 63262
rect 23662 63186 23714 63198
rect 25902 63250 25954 63262
rect 25902 63186 25954 63198
rect 27246 63250 27298 63262
rect 27246 63186 27298 63198
rect 27694 63250 27746 63262
rect 27694 63186 27746 63198
rect 28814 63250 28866 63262
rect 28814 63186 28866 63198
rect 2382 63138 2434 63150
rect 2382 63074 2434 63086
rect 7870 63138 7922 63150
rect 7870 63074 7922 63086
rect 8654 63138 8706 63150
rect 8654 63074 8706 63086
rect 9214 63138 9266 63150
rect 12238 63138 12290 63150
rect 11330 63086 11342 63138
rect 11394 63086 11406 63138
rect 9214 63074 9266 63086
rect 12238 63074 12290 63086
rect 13806 63138 13858 63150
rect 21758 63138 21810 63150
rect 14354 63086 14366 63138
rect 14418 63086 14430 63138
rect 16706 63086 16718 63138
rect 16770 63086 16782 63138
rect 17490 63086 17502 63138
rect 17554 63086 17566 63138
rect 18610 63086 18622 63138
rect 18674 63086 18686 63138
rect 13806 63074 13858 63086
rect 21758 63074 21810 63086
rect 21870 63138 21922 63150
rect 24222 63138 24274 63150
rect 22306 63086 22318 63138
rect 22370 63086 22382 63138
rect 21870 63074 21922 63086
rect 24222 63074 24274 63086
rect 25230 63138 25282 63150
rect 29922 63086 29934 63138
rect 29986 63086 29998 63138
rect 25230 63074 25282 63086
rect 13694 63026 13746 63038
rect 19630 63026 19682 63038
rect 17602 62974 17614 63026
rect 17666 62974 17678 63026
rect 13694 62962 13746 62974
rect 19630 62962 19682 62974
rect 19742 63026 19794 63038
rect 19742 62962 19794 62974
rect 25118 63026 25170 63038
rect 25118 62962 25170 62974
rect 28478 63026 28530 63038
rect 28478 62962 28530 62974
rect 29598 63026 29650 63038
rect 29598 62962 29650 62974
rect 4958 62914 5010 62926
rect 4958 62850 5010 62862
rect 6078 62914 6130 62926
rect 6078 62850 6130 62862
rect 7310 62914 7362 62926
rect 7310 62850 7362 62862
rect 9326 62914 9378 62926
rect 9326 62850 9378 62862
rect 9550 62914 9602 62926
rect 9550 62850 9602 62862
rect 20862 62914 20914 62926
rect 20862 62850 20914 62862
rect 21982 62914 22034 62926
rect 21982 62850 22034 62862
rect 22094 62914 22146 62926
rect 22094 62850 22146 62862
rect 24334 62914 24386 62926
rect 24334 62850 24386 62862
rect 26350 62914 26402 62926
rect 26350 62850 26402 62862
rect 26798 62914 26850 62926
rect 26798 62850 26850 62862
rect 29710 62914 29762 62926
rect 29710 62850 29762 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 1934 62578 1986 62590
rect 1934 62514 1986 62526
rect 2382 62578 2434 62590
rect 2382 62514 2434 62526
rect 2718 62578 2770 62590
rect 2718 62514 2770 62526
rect 3278 62578 3330 62590
rect 3278 62514 3330 62526
rect 3614 62578 3666 62590
rect 3614 62514 3666 62526
rect 4510 62578 4562 62590
rect 4510 62514 4562 62526
rect 5518 62578 5570 62590
rect 5518 62514 5570 62526
rect 5966 62578 6018 62590
rect 5966 62514 6018 62526
rect 6414 62578 6466 62590
rect 6414 62514 6466 62526
rect 7198 62578 7250 62590
rect 7198 62514 7250 62526
rect 7758 62578 7810 62590
rect 7758 62514 7810 62526
rect 8542 62578 8594 62590
rect 8542 62514 8594 62526
rect 8990 62578 9042 62590
rect 8990 62514 9042 62526
rect 10782 62578 10834 62590
rect 13358 62578 13410 62590
rect 12226 62526 12238 62578
rect 12290 62526 12302 62578
rect 10782 62514 10834 62526
rect 13358 62514 13410 62526
rect 13470 62578 13522 62590
rect 13470 62514 13522 62526
rect 13694 62578 13746 62590
rect 13694 62514 13746 62526
rect 15038 62578 15090 62590
rect 15038 62514 15090 62526
rect 15262 62578 15314 62590
rect 15262 62514 15314 62526
rect 15822 62578 15874 62590
rect 15822 62514 15874 62526
rect 16494 62578 16546 62590
rect 16494 62514 16546 62526
rect 16718 62578 16770 62590
rect 16718 62514 16770 62526
rect 19742 62578 19794 62590
rect 19742 62514 19794 62526
rect 20190 62578 20242 62590
rect 20190 62514 20242 62526
rect 20638 62578 20690 62590
rect 20638 62514 20690 62526
rect 21086 62578 21138 62590
rect 21086 62514 21138 62526
rect 21534 62578 21586 62590
rect 21534 62514 21586 62526
rect 22766 62578 22818 62590
rect 22766 62514 22818 62526
rect 23326 62578 23378 62590
rect 23326 62514 23378 62526
rect 23774 62578 23826 62590
rect 23774 62514 23826 62526
rect 24334 62578 24386 62590
rect 24334 62514 24386 62526
rect 24670 62578 24722 62590
rect 24670 62514 24722 62526
rect 25566 62578 25618 62590
rect 25566 62514 25618 62526
rect 26126 62578 26178 62590
rect 26126 62514 26178 62526
rect 26686 62578 26738 62590
rect 26686 62514 26738 62526
rect 27582 62578 27634 62590
rect 27582 62514 27634 62526
rect 28254 62578 28306 62590
rect 28254 62514 28306 62526
rect 28814 62578 28866 62590
rect 28814 62514 28866 62526
rect 11678 62466 11730 62478
rect 11678 62402 11730 62414
rect 15934 62466 15986 62478
rect 15934 62402 15986 62414
rect 22094 62466 22146 62478
rect 22094 62402 22146 62414
rect 22206 62466 22258 62478
rect 22206 62402 22258 62414
rect 28366 62466 28418 62478
rect 28366 62402 28418 62414
rect 4958 62354 5010 62366
rect 4834 62302 4846 62354
rect 4898 62302 4910 62354
rect 4174 62242 4226 62254
rect 4174 62178 4226 62190
rect 4849 62127 4895 62302
rect 4958 62290 5010 62302
rect 8094 62354 8146 62366
rect 8094 62290 8146 62302
rect 10558 62354 10610 62366
rect 10558 62290 10610 62302
rect 11230 62354 11282 62366
rect 11230 62290 11282 62302
rect 11902 62354 11954 62366
rect 11902 62290 11954 62302
rect 13582 62354 13634 62366
rect 14926 62354 14978 62366
rect 13906 62302 13918 62354
rect 13970 62302 13982 62354
rect 13582 62290 13634 62302
rect 14926 62290 14978 62302
rect 16830 62354 16882 62366
rect 16830 62290 16882 62302
rect 28030 62354 28082 62366
rect 28030 62290 28082 62302
rect 6750 62242 6802 62254
rect 6750 62178 6802 62190
rect 9998 62242 10050 62254
rect 9998 62178 10050 62190
rect 10670 62242 10722 62254
rect 10670 62178 10722 62190
rect 12686 62242 12738 62254
rect 12686 62178 12738 62190
rect 14366 62242 14418 62254
rect 14366 62178 14418 62190
rect 17950 62242 18002 62254
rect 17950 62178 18002 62190
rect 19294 62242 19346 62254
rect 19294 62178 19346 62190
rect 15710 62130 15762 62142
rect 8418 62127 8430 62130
rect 4849 62081 8430 62127
rect 8418 62078 8430 62081
rect 8482 62078 8494 62130
rect 12450 62078 12462 62130
rect 12514 62127 12526 62130
rect 12674 62127 12686 62130
rect 12514 62081 12686 62127
rect 12514 62078 12526 62081
rect 12674 62078 12686 62081
rect 12738 62078 12750 62130
rect 15710 62066 15762 62078
rect 18174 62130 18226 62142
rect 18498 62078 18510 62130
rect 18562 62078 18574 62130
rect 18174 62066 18226 62078
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 12574 61794 12626 61806
rect 3378 61742 3390 61794
rect 3442 61791 3454 61794
rect 4050 61791 4062 61794
rect 3442 61745 4062 61791
rect 3442 61742 3454 61745
rect 4050 61742 4062 61745
rect 4114 61742 4126 61794
rect 6290 61742 6302 61794
rect 6354 61791 6366 61794
rect 6738 61791 6750 61794
rect 6354 61745 6750 61791
rect 6354 61742 6366 61745
rect 6738 61742 6750 61745
rect 6802 61791 6814 61794
rect 7410 61791 7422 61794
rect 6802 61745 7422 61791
rect 6802 61742 6814 61745
rect 7410 61742 7422 61745
rect 7474 61742 7486 61794
rect 12574 61730 12626 61742
rect 12910 61794 12962 61806
rect 12910 61730 12962 61742
rect 15710 61794 15762 61806
rect 15710 61730 15762 61742
rect 16158 61794 16210 61806
rect 17266 61742 17278 61794
rect 17330 61791 17342 61794
rect 17490 61791 17502 61794
rect 17330 61745 17502 61791
rect 17330 61742 17342 61745
rect 17490 61742 17502 61745
rect 17554 61791 17566 61794
rect 17938 61791 17950 61794
rect 17554 61745 17950 61791
rect 17554 61742 17566 61745
rect 17938 61742 17950 61745
rect 18002 61742 18014 61794
rect 21858 61742 21870 61794
rect 21922 61791 21934 61794
rect 22418 61791 22430 61794
rect 21922 61745 22430 61791
rect 21922 61742 21934 61745
rect 22418 61742 22430 61745
rect 22482 61742 22494 61794
rect 16158 61730 16210 61742
rect 2382 61682 2434 61694
rect 2382 61618 2434 61630
rect 2718 61682 2770 61694
rect 2718 61618 2770 61630
rect 3166 61682 3218 61694
rect 3166 61618 3218 61630
rect 4510 61682 4562 61694
rect 4510 61618 4562 61630
rect 4958 61682 5010 61694
rect 4958 61618 5010 61630
rect 5854 61682 5906 61694
rect 5854 61618 5906 61630
rect 6302 61682 6354 61694
rect 6302 61618 6354 61630
rect 7198 61682 7250 61694
rect 7198 61618 7250 61630
rect 7758 61682 7810 61694
rect 7758 61618 7810 61630
rect 8878 61682 8930 61694
rect 8878 61618 8930 61630
rect 9326 61682 9378 61694
rect 9326 61618 9378 61630
rect 9886 61682 9938 61694
rect 9886 61618 9938 61630
rect 10782 61682 10834 61694
rect 10782 61618 10834 61630
rect 10894 61682 10946 61694
rect 10894 61618 10946 61630
rect 11566 61682 11618 61694
rect 11566 61618 11618 61630
rect 13806 61682 13858 61694
rect 13806 61618 13858 61630
rect 17166 61682 17218 61694
rect 17166 61618 17218 61630
rect 20750 61682 20802 61694
rect 20750 61618 20802 61630
rect 21758 61682 21810 61694
rect 21758 61618 21810 61630
rect 22206 61682 22258 61694
rect 22206 61618 22258 61630
rect 23550 61682 23602 61694
rect 23550 61618 23602 61630
rect 24222 61682 24274 61694
rect 24222 61618 24274 61630
rect 25006 61682 25058 61694
rect 25006 61618 25058 61630
rect 25342 61682 25394 61694
rect 25342 61618 25394 61630
rect 25902 61682 25954 61694
rect 25902 61618 25954 61630
rect 4062 61570 4114 61582
rect 4062 61506 4114 61518
rect 6750 61570 6802 61582
rect 6750 61506 6802 61518
rect 10222 61570 10274 61582
rect 14366 61570 14418 61582
rect 11106 61518 11118 61570
rect 11170 61518 11182 61570
rect 12562 61518 12574 61570
rect 12626 61518 12638 61570
rect 10222 61506 10274 61518
rect 14366 61506 14418 61518
rect 15150 61570 15202 61582
rect 15150 61506 15202 61518
rect 15822 61570 15874 61582
rect 15822 61506 15874 61518
rect 16046 61570 16098 61582
rect 16046 61506 16098 61518
rect 19742 61570 19794 61582
rect 19742 61506 19794 61518
rect 14702 61458 14754 61470
rect 14702 61394 14754 61406
rect 16718 61458 16770 61470
rect 16718 61394 16770 61406
rect 1934 61346 1986 61358
rect 1934 61282 1986 61294
rect 3614 61346 3666 61358
rect 3614 61282 3666 61294
rect 8430 61346 8482 61358
rect 8430 61282 8482 61294
rect 12014 61346 12066 61358
rect 12014 61282 12066 61294
rect 13694 61346 13746 61358
rect 13694 61282 13746 61294
rect 13918 61346 13970 61358
rect 13918 61282 13970 61294
rect 17614 61346 17666 61358
rect 17614 61282 17666 61294
rect 18062 61346 18114 61358
rect 18062 61282 18114 61294
rect 18734 61346 18786 61358
rect 18734 61282 18786 61294
rect 19182 61346 19234 61358
rect 19182 61282 19234 61294
rect 20302 61346 20354 61358
rect 20302 61282 20354 61294
rect 22654 61346 22706 61358
rect 22654 61282 22706 61294
rect 23102 61346 23154 61358
rect 23102 61282 23154 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 1934 61010 1986 61022
rect 1934 60946 1986 60958
rect 2382 61010 2434 61022
rect 2382 60946 2434 60958
rect 2830 61010 2882 61022
rect 2830 60946 2882 60958
rect 3166 61010 3218 61022
rect 3166 60946 3218 60958
rect 4174 61010 4226 61022
rect 4174 60946 4226 60958
rect 4958 61010 5010 61022
rect 4958 60946 5010 60958
rect 5854 61010 5906 61022
rect 5854 60946 5906 60958
rect 6862 61010 6914 61022
rect 6862 60946 6914 60958
rect 8654 61010 8706 61022
rect 8654 60946 8706 60958
rect 10110 61010 10162 61022
rect 10110 60946 10162 60958
rect 10222 61010 10274 61022
rect 10222 60946 10274 60958
rect 10782 61010 10834 61022
rect 10782 60946 10834 60958
rect 13470 61010 13522 61022
rect 13470 60946 13522 60958
rect 13694 61010 13746 61022
rect 13694 60946 13746 60958
rect 14478 61010 14530 61022
rect 14478 60946 14530 60958
rect 15038 61010 15090 61022
rect 15038 60946 15090 60958
rect 15374 61010 15426 61022
rect 15374 60946 15426 60958
rect 17054 61010 17106 61022
rect 17054 60946 17106 60958
rect 18286 61010 18338 61022
rect 18286 60946 18338 60958
rect 19742 61010 19794 61022
rect 19742 60946 19794 60958
rect 20638 61010 20690 61022
rect 20638 60946 20690 60958
rect 21870 61010 21922 61022
rect 21870 60946 21922 60958
rect 22318 61010 22370 61022
rect 22318 60946 22370 60958
rect 22654 61010 22706 61022
rect 22654 60946 22706 60958
rect 23550 61010 23602 61022
rect 23550 60946 23602 60958
rect 24110 61010 24162 61022
rect 24110 60946 24162 60958
rect 29822 61010 29874 61022
rect 29822 60946 29874 60958
rect 30382 61010 30434 61022
rect 30382 60946 30434 60958
rect 30942 61010 30994 61022
rect 30942 60946 30994 60958
rect 7758 60898 7810 60910
rect 7758 60834 7810 60846
rect 13358 60898 13410 60910
rect 13358 60834 13410 60846
rect 14030 60898 14082 60910
rect 14030 60834 14082 60846
rect 15822 60898 15874 60910
rect 15822 60834 15874 60846
rect 17614 60898 17666 60910
rect 17614 60834 17666 60846
rect 30270 60898 30322 60910
rect 30270 60834 30322 60846
rect 5518 60786 5570 60798
rect 5518 60722 5570 60734
rect 6302 60786 6354 60798
rect 6302 60722 6354 60734
rect 19182 60786 19234 60798
rect 19182 60722 19234 60734
rect 3726 60674 3778 60686
rect 3726 60610 3778 60622
rect 4510 60674 4562 60686
rect 4510 60610 4562 60622
rect 7198 60674 7250 60686
rect 7198 60610 7250 60622
rect 8094 60674 8146 60686
rect 8094 60610 8146 60622
rect 8990 60674 9042 60686
rect 8990 60610 9042 60622
rect 11454 60674 11506 60686
rect 11454 60610 11506 60622
rect 11902 60674 11954 60686
rect 11902 60610 11954 60622
rect 12350 60674 12402 60686
rect 12350 60610 12402 60622
rect 12798 60674 12850 60686
rect 12798 60610 12850 60622
rect 16270 60674 16322 60686
rect 16270 60610 16322 60622
rect 18734 60674 18786 60686
rect 18734 60610 18786 60622
rect 20190 60674 20242 60686
rect 20190 60610 20242 60622
rect 21310 60674 21362 60686
rect 21310 60610 21362 60622
rect 23214 60674 23266 60686
rect 23214 60610 23266 60622
rect 9998 60562 10050 60574
rect 30382 60562 30434 60574
rect 18722 60510 18734 60562
rect 18786 60559 18798 60562
rect 19394 60559 19406 60562
rect 18786 60513 19406 60559
rect 18786 60510 18798 60513
rect 19394 60510 19406 60513
rect 19458 60510 19470 60562
rect 9998 60498 10050 60510
rect 30382 60498 30434 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 3490 60174 3502 60226
rect 3554 60223 3566 60226
rect 4834 60223 4846 60226
rect 3554 60177 4846 60223
rect 3554 60174 3566 60177
rect 4834 60174 4846 60177
rect 4898 60174 4910 60226
rect 2158 60114 2210 60126
rect 2158 60050 2210 60062
rect 2606 60114 2658 60126
rect 2606 60050 2658 60062
rect 3054 60114 3106 60126
rect 3054 60050 3106 60062
rect 3390 60114 3442 60126
rect 3390 60050 3442 60062
rect 3950 60114 4002 60126
rect 3950 60050 4002 60062
rect 4846 60114 4898 60126
rect 4846 60050 4898 60062
rect 7758 60114 7810 60126
rect 7758 60050 7810 60062
rect 8206 60114 8258 60126
rect 8206 60050 8258 60062
rect 8654 60114 8706 60126
rect 8654 60050 8706 60062
rect 8990 60114 9042 60126
rect 8990 60050 9042 60062
rect 9438 60114 9490 60126
rect 9438 60050 9490 60062
rect 10670 60114 10722 60126
rect 10670 60050 10722 60062
rect 11230 60114 11282 60126
rect 13582 60114 13634 60126
rect 12674 60062 12686 60114
rect 12738 60062 12750 60114
rect 11230 60050 11282 60062
rect 13582 60050 13634 60062
rect 14254 60114 14306 60126
rect 14254 60050 14306 60062
rect 14702 60114 14754 60126
rect 14702 60050 14754 60062
rect 15822 60114 15874 60126
rect 15822 60050 15874 60062
rect 16382 60114 16434 60126
rect 16382 60050 16434 60062
rect 16830 60114 16882 60126
rect 16830 60050 16882 60062
rect 17614 60114 17666 60126
rect 17614 60050 17666 60062
rect 19518 60114 19570 60126
rect 19518 60050 19570 60062
rect 20414 60114 20466 60126
rect 20414 60050 20466 60062
rect 20862 60114 20914 60126
rect 20862 60050 20914 60062
rect 21982 60114 22034 60126
rect 21982 60050 22034 60062
rect 23214 60114 23266 60126
rect 23214 60050 23266 60062
rect 23662 60114 23714 60126
rect 23662 60050 23714 60062
rect 6302 60002 6354 60014
rect 18286 60002 18338 60014
rect 11666 59950 11678 60002
rect 11730 59950 11742 60002
rect 6302 59938 6354 59950
rect 18286 59938 18338 59950
rect 9998 59890 10050 59902
rect 9998 59826 10050 59838
rect 15374 59890 15426 59902
rect 15374 59826 15426 59838
rect 19070 59890 19122 59902
rect 19070 59826 19122 59838
rect 4398 59778 4450 59790
rect 4398 59714 4450 59726
rect 5854 59778 5906 59790
rect 5854 59714 5906 59726
rect 6638 59778 6690 59790
rect 6638 59714 6690 59726
rect 7086 59778 7138 59790
rect 7086 59714 7138 59726
rect 17278 59778 17330 59790
rect 17278 59714 17330 59726
rect 19854 59778 19906 59790
rect 19854 59714 19906 59726
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 3950 59442 4002 59454
rect 3950 59378 4002 59390
rect 4734 59442 4786 59454
rect 4734 59378 4786 59390
rect 5294 59442 5346 59454
rect 5294 59378 5346 59390
rect 6302 59442 6354 59454
rect 6302 59378 6354 59390
rect 6862 59442 6914 59454
rect 6862 59378 6914 59390
rect 7310 59442 7362 59454
rect 7310 59378 7362 59390
rect 8654 59442 8706 59454
rect 8654 59378 8706 59390
rect 9102 59442 9154 59454
rect 9102 59378 9154 59390
rect 9774 59442 9826 59454
rect 9774 59378 9826 59390
rect 11230 59442 11282 59454
rect 11230 59378 11282 59390
rect 11678 59442 11730 59454
rect 11678 59378 11730 59390
rect 12462 59442 12514 59454
rect 12462 59378 12514 59390
rect 13022 59442 13074 59454
rect 13022 59378 13074 59390
rect 14926 59442 14978 59454
rect 14926 59378 14978 59390
rect 15486 59442 15538 59454
rect 15486 59378 15538 59390
rect 15934 59442 15986 59454
rect 15934 59378 15986 59390
rect 16494 59442 16546 59454
rect 16494 59378 16546 59390
rect 16942 59442 16994 59454
rect 16942 59378 16994 59390
rect 17726 59442 17778 59454
rect 17726 59378 17778 59390
rect 18510 59442 18562 59454
rect 18510 59378 18562 59390
rect 13582 59330 13634 59342
rect 13582 59266 13634 59278
rect 3390 59106 3442 59118
rect 3390 59042 3442 59054
rect 4398 59106 4450 59118
rect 4398 59042 4450 59054
rect 5966 59106 6018 59118
rect 5966 59042 6018 59054
rect 7646 59106 7698 59118
rect 7646 59042 7698 59054
rect 8094 59106 8146 59118
rect 8094 59042 8146 59054
rect 10446 59106 10498 59118
rect 10446 59042 10498 59054
rect 10782 59106 10834 59118
rect 10782 59042 10834 59054
rect 14030 59106 14082 59118
rect 14030 59042 14082 59054
rect 18174 59106 18226 59118
rect 18174 59042 18226 59054
rect 18958 59106 19010 59118
rect 18958 59042 19010 59054
rect 6066 58942 6078 58994
rect 6130 58991 6142 58994
rect 6626 58991 6638 58994
rect 6130 58945 6638 58991
rect 6130 58942 6142 58945
rect 6626 58942 6638 58945
rect 6690 58942 6702 58994
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 19518 58658 19570 58670
rect 15586 58606 15598 58658
rect 15650 58655 15662 58658
rect 16258 58655 16270 58658
rect 15650 58609 16270 58655
rect 15650 58606 15662 58609
rect 16258 58606 16270 58609
rect 16322 58606 16334 58658
rect 19518 58594 19570 58606
rect 4062 58546 4114 58558
rect 4062 58482 4114 58494
rect 5854 58546 5906 58558
rect 5854 58482 5906 58494
rect 6302 58546 6354 58558
rect 6302 58482 6354 58494
rect 9326 58546 9378 58558
rect 9326 58482 9378 58494
rect 9774 58546 9826 58558
rect 9774 58482 9826 58494
rect 10222 58546 10274 58558
rect 10222 58482 10274 58494
rect 11230 58546 11282 58558
rect 11230 58482 11282 58494
rect 11678 58546 11730 58558
rect 11678 58482 11730 58494
rect 12126 58546 12178 58558
rect 12126 58482 12178 58494
rect 12574 58546 12626 58558
rect 12574 58482 12626 58494
rect 13022 58546 13074 58558
rect 13022 58482 13074 58494
rect 13694 58546 13746 58558
rect 13694 58482 13746 58494
rect 15038 58546 15090 58558
rect 15038 58482 15090 58494
rect 15374 58546 15426 58558
rect 15374 58482 15426 58494
rect 15934 58546 15986 58558
rect 15934 58482 15986 58494
rect 16270 58546 16322 58558
rect 16270 58482 16322 58494
rect 17166 58546 17218 58558
rect 17166 58482 17218 58494
rect 17726 58546 17778 58558
rect 17726 58482 17778 58494
rect 18174 58546 18226 58558
rect 18174 58482 18226 58494
rect 19630 58546 19682 58558
rect 19630 58482 19682 58494
rect 20078 58546 20130 58558
rect 20078 58482 20130 58494
rect 10670 58434 10722 58446
rect 10670 58370 10722 58382
rect 6750 58210 6802 58222
rect 6750 58146 6802 58158
rect 7198 58210 7250 58222
rect 7198 58146 7250 58158
rect 7646 58210 7698 58222
rect 7646 58146 7698 58158
rect 8094 58210 8146 58222
rect 8094 58146 8146 58158
rect 8766 58210 8818 58222
rect 8766 58146 8818 58158
rect 14030 58210 14082 58222
rect 14030 58146 14082 58158
rect 14478 58210 14530 58222
rect 14478 58146 14530 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 7870 57874 7922 57886
rect 7870 57810 7922 57822
rect 8318 57874 8370 57886
rect 8318 57810 8370 57822
rect 8990 57874 9042 57886
rect 8990 57810 9042 57822
rect 9774 57874 9826 57886
rect 9774 57810 9826 57822
rect 10446 57874 10498 57886
rect 10446 57810 10498 57822
rect 11118 57874 11170 57886
rect 11118 57810 11170 57822
rect 11566 57874 11618 57886
rect 11566 57810 11618 57822
rect 12014 57874 12066 57886
rect 12014 57810 12066 57822
rect 12462 57874 12514 57886
rect 12462 57810 12514 57822
rect 13022 57874 13074 57886
rect 13022 57810 13074 57822
rect 15150 57874 15202 57886
rect 15150 57810 15202 57822
rect 13806 57762 13858 57774
rect 13806 57698 13858 57710
rect 14254 57650 14306 57662
rect 14254 57586 14306 57598
rect 7310 57538 7362 57550
rect 7310 57474 7362 57486
rect 13358 57538 13410 57550
rect 13358 57474 13410 57486
rect 14702 57538 14754 57550
rect 14702 57474 14754 57486
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 9326 56978 9378 56990
rect 9326 56914 9378 56926
rect 9774 56978 9826 56990
rect 9774 56914 9826 56926
rect 10222 56978 10274 56990
rect 10222 56914 10274 56926
rect 14142 56978 14194 56990
rect 14142 56914 14194 56926
rect 13582 56866 13634 56878
rect 13582 56802 13634 56814
rect 12574 56642 12626 56654
rect 12574 56578 12626 56590
rect 12910 56642 12962 56654
rect 12910 56578 12962 56590
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 28814 55298 28866 55310
rect 28814 55234 28866 55246
rect 29598 55298 29650 55310
rect 29598 55234 29650 55246
rect 29934 55074 29986 55086
rect 29934 55010 29986 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 17614 36706 17666 36718
rect 17614 36642 17666 36654
rect 16942 36594 16994 36606
rect 16942 36530 16994 36542
rect 17490 36430 17502 36482
rect 17554 36430 17566 36482
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 12462 6130 12514 6142
rect 12462 6066 12514 6078
rect 14366 6130 14418 6142
rect 14366 6066 14418 6078
rect 14814 6130 14866 6142
rect 14814 6066 14866 6078
rect 51214 6130 51266 6142
rect 51214 6066 51266 6078
rect 19630 6018 19682 6030
rect 19630 5954 19682 5966
rect 11006 5906 11058 5918
rect 11006 5842 11058 5854
rect 18622 5906 18674 5918
rect 18622 5842 18674 5854
rect 52222 5906 52274 5918
rect 52222 5842 52274 5854
rect 12126 5794 12178 5806
rect 12126 5730 12178 5742
rect 15374 5794 15426 5806
rect 15374 5730 15426 5742
rect 18174 5794 18226 5806
rect 18174 5730 18226 5742
rect 34302 5794 34354 5806
rect 34302 5730 34354 5742
rect 51774 5794 51826 5806
rect 51774 5730 51826 5742
rect 11230 5682 11282 5694
rect 18846 5682 18898 5694
rect 52446 5682 52498 5694
rect 11554 5630 11566 5682
rect 11618 5630 11630 5682
rect 19170 5630 19182 5682
rect 19234 5630 19246 5682
rect 52770 5630 52782 5682
rect 52834 5630 52846 5682
rect 11230 5618 11282 5630
rect 18846 5618 18898 5630
rect 52446 5618 52498 5630
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 22766 5234 22818 5246
rect 22766 5170 22818 5182
rect 23214 5234 23266 5246
rect 23214 5170 23266 5182
rect 32622 5234 32674 5246
rect 32622 5170 32674 5182
rect 33070 5234 33122 5246
rect 33070 5170 33122 5182
rect 34302 5234 34354 5246
rect 34302 5170 34354 5182
rect 34750 5234 34802 5246
rect 34750 5170 34802 5182
rect 40014 5234 40066 5246
rect 40014 5170 40066 5182
rect 40462 5234 40514 5246
rect 40462 5170 40514 5182
rect 46846 5234 46898 5246
rect 46846 5170 46898 5182
rect 47742 5234 47794 5246
rect 47742 5170 47794 5182
rect 53342 5234 53394 5246
rect 53342 5170 53394 5182
rect 22206 5122 22258 5134
rect 11442 5070 11454 5122
rect 11506 5070 11518 5122
rect 22206 5058 22258 5070
rect 23438 5122 23490 5134
rect 23438 5058 23490 5070
rect 32062 5122 32114 5134
rect 32062 5058 32114 5070
rect 33294 5122 33346 5134
rect 33294 5058 33346 5070
rect 34974 5122 35026 5134
rect 34974 5058 35026 5070
rect 39454 5122 39506 5134
rect 39454 5058 39506 5070
rect 40686 5122 40738 5134
rect 40686 5058 40738 5070
rect 47182 5122 47234 5134
rect 47182 5058 47234 5070
rect 47966 5122 48018 5134
rect 47966 5058 48018 5070
rect 52334 5122 52386 5134
rect 52334 5058 52386 5070
rect 24334 5010 24386 5022
rect 23762 4958 23774 5010
rect 23826 4958 23838 5010
rect 24334 4946 24386 4958
rect 11678 4898 11730 4910
rect 11678 4834 11730 4846
rect 24670 4898 24722 4910
rect 33618 4846 33630 4898
rect 33682 4846 33694 4898
rect 35298 4846 35310 4898
rect 35362 4846 35374 4898
rect 41010 4846 41022 4898
rect 41074 4846 41086 4898
rect 48290 4846 48302 4898
rect 48354 4846 48366 4898
rect 24670 4834 24722 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 12350 4562 12402 4574
rect 12350 4498 12402 4510
rect 14590 4562 14642 4574
rect 14590 4498 14642 4510
rect 26798 4562 26850 4574
rect 26798 4498 26850 4510
rect 27246 4562 27298 4574
rect 27246 4498 27298 4510
rect 50766 4562 50818 4574
rect 50766 4498 50818 4510
rect 51214 4562 51266 4574
rect 51214 4498 51266 4510
rect 7310 4450 7362 4462
rect 7310 4386 7362 4398
rect 12798 4450 12850 4462
rect 12798 4386 12850 4398
rect 16606 4450 16658 4462
rect 16606 4386 16658 4398
rect 19630 4450 19682 4462
rect 19630 4386 19682 4398
rect 19966 4450 20018 4462
rect 19966 4386 20018 4398
rect 29598 4450 29650 4462
rect 29598 4386 29650 4398
rect 34302 4450 34354 4462
rect 34302 4386 34354 4398
rect 34638 4450 34690 4462
rect 34638 4386 34690 4398
rect 38334 4450 38386 4462
rect 38334 4386 38386 4398
rect 38670 4450 38722 4462
rect 38670 4386 38722 4398
rect 43486 4450 43538 4462
rect 43486 4386 43538 4398
rect 43822 4450 43874 4462
rect 43822 4386 43874 4398
rect 49534 4450 49586 4462
rect 49534 4386 49586 4398
rect 49870 4450 49922 4462
rect 49870 4386 49922 4398
rect 54350 4450 54402 4462
rect 54350 4386 54402 4398
rect 54910 4450 54962 4462
rect 54910 4386 54962 4398
rect 55246 4450 55298 4462
rect 55246 4386 55298 4398
rect 58270 4450 58322 4462
rect 58270 4386 58322 4398
rect 66222 4450 66274 4462
rect 66222 4386 66274 4398
rect 7646 4338 7698 4350
rect 11678 4338 11730 4350
rect 11330 4286 11342 4338
rect 11394 4286 11406 4338
rect 7646 4274 7698 4286
rect 11678 4274 11730 4286
rect 11902 4338 11954 4350
rect 11902 4274 11954 4286
rect 15150 4338 15202 4350
rect 15150 4274 15202 4286
rect 15374 4338 15426 4350
rect 16270 4338 16322 4350
rect 15698 4286 15710 4338
rect 15762 4286 15774 4338
rect 15374 4274 15426 4286
rect 16270 4274 16322 4286
rect 27806 4338 27858 4350
rect 27806 4274 27858 4286
rect 28030 4338 28082 4350
rect 29262 4338 29314 4350
rect 28354 4286 28366 4338
rect 28418 4286 28430 4338
rect 28030 4274 28082 4286
rect 29262 4274 29314 4286
rect 51774 4338 51826 4350
rect 51774 4274 51826 4286
rect 51998 4338 52050 4350
rect 51998 4274 52050 4286
rect 52894 4338 52946 4350
rect 52894 4274 52946 4286
rect 53118 4338 53170 4350
rect 54014 4338 54066 4350
rect 53442 4286 53454 4338
rect 53506 4286 53518 4338
rect 53118 4274 53170 4286
rect 54014 4274 54066 4286
rect 57934 4338 57986 4350
rect 57934 4274 57986 4286
rect 65886 4338 65938 4350
rect 65886 4274 65938 4286
rect 74398 4338 74450 4350
rect 75170 4286 75182 4338
rect 75234 4286 75246 4338
rect 74398 4274 74450 4286
rect 65326 4226 65378 4238
rect 52322 4174 52334 4226
rect 52386 4174 52398 4226
rect 76066 4174 76078 4226
rect 76130 4174 76142 4226
rect 65326 4162 65378 4174
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 53006 3778 53058 3790
rect 53006 3714 53058 3726
rect 16046 3666 16098 3678
rect 52110 3666 52162 3678
rect 7858 3614 7870 3666
rect 7922 3614 7934 3666
rect 12226 3614 12238 3666
rect 12290 3614 12302 3666
rect 18162 3614 18174 3666
rect 18226 3614 18238 3666
rect 22082 3614 22094 3666
rect 22146 3614 22158 3666
rect 26674 3614 26686 3666
rect 26738 3614 26750 3666
rect 31378 3614 31390 3666
rect 31442 3614 31454 3666
rect 35746 3614 35758 3666
rect 35810 3614 35822 3666
rect 41682 3614 41694 3666
rect 41746 3614 41758 3666
rect 45602 3614 45614 3666
rect 45666 3614 45678 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 59266 3614 59278 3666
rect 59330 3614 59342 3666
rect 65202 3614 65214 3666
rect 65266 3614 65278 3666
rect 69122 3614 69134 3666
rect 69186 3614 69198 3666
rect 73714 3614 73726 3666
rect 73778 3614 73790 3666
rect 16046 3602 16098 3614
rect 52110 3602 52162 3614
rect 4286 3554 4338 3566
rect 51662 3554 51714 3566
rect 3490 3502 3502 3554
rect 3554 3502 3566 3554
rect 7298 3502 7310 3554
rect 7362 3502 7374 3554
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 17490 3502 17502 3554
rect 17554 3502 17566 3554
rect 21410 3502 21422 3554
rect 21474 3502 21486 3554
rect 26002 3502 26014 3554
rect 26066 3502 26078 3554
rect 30706 3502 30718 3554
rect 30770 3502 30782 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 41010 3502 41022 3554
rect 41074 3502 41086 3554
rect 44930 3502 44942 3554
rect 44994 3502 45006 3554
rect 50530 3502 50542 3554
rect 50594 3502 50606 3554
rect 4286 3490 4338 3502
rect 51662 3490 51714 3502
rect 52782 3554 52834 3566
rect 72606 3554 72658 3566
rect 53330 3502 53342 3554
rect 53394 3502 53406 3554
rect 54338 3502 54350 3554
rect 54402 3502 54414 3554
rect 58594 3502 58606 3554
rect 58658 3502 58670 3554
rect 64530 3502 64542 3554
rect 64594 3502 64606 3554
rect 68450 3502 68462 3554
rect 68514 3502 68526 3554
rect 73266 3502 73278 3554
rect 73330 3502 73342 3554
rect 52782 3490 52834 3502
rect 72606 3490 72658 3502
rect 2594 3390 2606 3442
rect 2658 3390 2670 3442
rect 49634 3390 49646 3442
rect 49698 3390 49710 3442
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
<< via1 >>
rect 7086 77646 7138 77698
rect 9662 77646 9714 77698
rect 11790 76974 11842 77026
rect 12350 76974 12402 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 2046 76638 2098 76690
rect 2494 76638 2546 76690
rect 2942 76638 2994 76690
rect 4734 76638 4786 76690
rect 5854 76638 5906 76690
rect 9998 76638 10050 76690
rect 37550 76638 37602 76690
rect 39902 76638 39954 76690
rect 40910 76638 40962 76690
rect 41918 76638 41970 76690
rect 59950 76638 60002 76690
rect 63870 76638 63922 76690
rect 67790 76638 67842 76690
rect 72494 76638 72546 76690
rect 3502 76526 3554 76578
rect 7534 76526 7586 76578
rect 12350 76526 12402 76578
rect 23550 76526 23602 76578
rect 27470 76526 27522 76578
rect 30606 76526 30658 76578
rect 31726 76526 31778 76578
rect 31838 76526 31890 76578
rect 34638 76526 34690 76578
rect 35982 76526 36034 76578
rect 39006 76526 39058 76578
rect 43374 76526 43426 76578
rect 47630 76526 47682 76578
rect 48750 76526 48802 76578
rect 51550 76526 51602 76578
rect 52670 76526 52722 76578
rect 61630 76526 61682 76578
rect 65550 76526 65602 76578
rect 69582 76526 69634 76578
rect 73950 76526 74002 76578
rect 3614 76414 3666 76466
rect 4398 76414 4450 76466
rect 4734 76414 4786 76466
rect 6302 76414 6354 76466
rect 6638 76414 6690 76466
rect 6862 76414 6914 76466
rect 10446 76414 10498 76466
rect 10558 76414 10610 76466
rect 10670 76414 10722 76466
rect 16718 76414 16770 76466
rect 17726 76414 17778 76466
rect 24334 76414 24386 76466
rect 28142 76414 28194 76466
rect 32062 76414 32114 76466
rect 6750 76302 6802 76354
rect 8878 76302 8930 76354
rect 11566 76302 11618 76354
rect 13806 76302 13858 76354
rect 15934 76302 15986 76354
rect 18510 76302 18562 76354
rect 20638 76302 20690 76354
rect 21422 76302 21474 76354
rect 25342 76302 25394 76354
rect 29486 76302 29538 76354
rect 33182 76302 33234 76354
rect 33630 76302 33682 76354
rect 35646 76302 35698 76354
rect 37102 76302 37154 76354
rect 37998 76302 38050 76354
rect 41358 76302 41410 76354
rect 42366 76302 42418 76354
rect 46622 76302 46674 76354
rect 50542 76302 50594 76354
rect 60622 76302 60674 76354
rect 64542 76302 64594 76354
rect 68574 76302 68626 76354
rect 72942 76302 72994 76354
rect 3726 76190 3778 76242
rect 4622 76190 4674 76242
rect 31278 76190 31330 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 2046 75854 2098 75906
rect 37326 75854 37378 75906
rect 37998 75854 38050 75906
rect 3614 75742 3666 75794
rect 6078 75742 6130 75794
rect 8206 75742 8258 75794
rect 12910 75742 12962 75794
rect 14590 75742 14642 75794
rect 16830 75742 16882 75794
rect 19406 75742 19458 75794
rect 22990 75742 23042 75794
rect 25118 75742 25170 75794
rect 28030 75742 28082 75794
rect 29822 75742 29874 75794
rect 31054 75742 31106 75794
rect 36542 75742 36594 75794
rect 4062 75686 4114 75738
rect 38334 75742 38386 75794
rect 38782 75742 38834 75794
rect 40126 75742 40178 75794
rect 55022 75742 55074 75794
rect 55470 75742 55522 75794
rect 74958 75742 75010 75794
rect 77198 75742 77250 75794
rect 4286 75630 4338 75682
rect 4510 75630 4562 75682
rect 8990 75630 9042 75682
rect 10110 75630 10162 75682
rect 13582 75630 13634 75682
rect 17502 75630 17554 75682
rect 21758 75630 21810 75682
rect 22318 75630 22370 75682
rect 28702 75630 28754 75682
rect 30942 75630 30994 75682
rect 31950 75630 32002 75682
rect 32398 75630 32450 75682
rect 32846 75630 32898 75682
rect 34190 75630 34242 75682
rect 34974 75630 35026 75682
rect 4734 75518 4786 75570
rect 4958 75518 5010 75570
rect 10782 75518 10834 75570
rect 13918 75518 13970 75570
rect 18622 75518 18674 75570
rect 20414 75518 20466 75570
rect 31390 75518 31442 75570
rect 32958 75518 33010 75570
rect 33406 75518 33458 75570
rect 36094 75518 36146 75570
rect 56478 75518 56530 75570
rect 76302 75518 76354 75570
rect 2830 75406 2882 75458
rect 4510 75406 4562 75458
rect 9550 75406 9602 75458
rect 13806 75406 13858 75458
rect 18174 75406 18226 75458
rect 18286 75406 18338 75458
rect 18398 75406 18450 75458
rect 25790 75406 25842 75458
rect 35758 75406 35810 75458
rect 37438 75406 37490 75458
rect 37886 75406 37938 75458
rect 39230 75406 39282 75458
rect 39678 75406 39730 75458
rect 40574 75406 40626 75458
rect 41022 75406 41074 75458
rect 41470 75406 41522 75458
rect 41918 75406 41970 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 2382 75070 2434 75122
rect 12350 75070 12402 75122
rect 35422 75070 35474 75122
rect 35870 75070 35922 75122
rect 38558 75070 38610 75122
rect 39454 75070 39506 75122
rect 7758 74958 7810 75010
rect 11342 74958 11394 75010
rect 13022 74958 13074 75010
rect 13134 74958 13186 75010
rect 18734 74958 18786 75010
rect 24894 74958 24946 75010
rect 27806 74958 27858 75010
rect 31838 74958 31890 75010
rect 33742 74958 33794 75010
rect 3166 74846 3218 74898
rect 6862 74846 6914 74898
rect 8430 74846 8482 74898
rect 8766 74846 8818 74898
rect 8990 74846 9042 74898
rect 11118 74846 11170 74898
rect 11454 74846 11506 74898
rect 12574 74846 12626 74898
rect 16942 74846 16994 74898
rect 20302 74846 20354 74898
rect 24222 74846 24274 74898
rect 24446 74846 24498 74898
rect 24670 74846 24722 74898
rect 28590 74846 28642 74898
rect 29710 74846 29762 74898
rect 30830 74846 30882 74898
rect 31166 74846 31218 74898
rect 31950 74846 32002 74898
rect 32398 74846 32450 74898
rect 34302 74846 34354 74898
rect 34526 74846 34578 74898
rect 1934 74734 1986 74786
rect 3838 74734 3890 74786
rect 6078 74734 6130 74786
rect 8542 74734 8594 74786
rect 10558 74734 10610 74786
rect 13358 74734 13410 74786
rect 14030 74734 14082 74786
rect 16158 74734 16210 74786
rect 17726 74734 17778 74786
rect 19854 74734 19906 74786
rect 21086 74734 21138 74786
rect 23214 74734 23266 74786
rect 25678 74734 25730 74786
rect 29038 74734 29090 74786
rect 32846 74734 32898 74786
rect 34974 74734 35026 74786
rect 36318 74734 36370 74786
rect 36766 74734 36818 74786
rect 37214 74734 37266 74786
rect 37662 74734 37714 74786
rect 38110 74734 38162 74786
rect 39006 74734 39058 74786
rect 39902 74734 39954 74786
rect 40350 74734 40402 74786
rect 40798 74734 40850 74786
rect 41470 74734 41522 74786
rect 2830 74622 2882 74674
rect 3166 74622 3218 74674
rect 7534 74622 7586 74674
rect 7870 74622 7922 74674
rect 9998 74622 10050 74674
rect 10334 74622 10386 74674
rect 11902 74622 11954 74674
rect 24782 74622 24834 74674
rect 33854 74622 33906 74674
rect 34078 74622 34130 74674
rect 37550 74622 37602 74674
rect 39006 74622 39058 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 2942 74286 2994 74338
rect 3278 74286 3330 74338
rect 7086 74286 7138 74338
rect 9662 74286 9714 74338
rect 11230 74286 11282 74338
rect 11790 74286 11842 74338
rect 37326 74286 37378 74338
rect 38110 74286 38162 74338
rect 38670 74286 38722 74338
rect 39902 74286 39954 74338
rect 2158 74174 2210 74226
rect 2606 74174 2658 74226
rect 3054 74174 3106 74226
rect 4846 74174 4898 74226
rect 5966 74174 6018 74226
rect 14478 74174 14530 74226
rect 16606 74174 16658 74226
rect 17950 74174 18002 74226
rect 20078 74174 20130 74226
rect 26350 74174 26402 74226
rect 27022 74174 27074 74226
rect 30606 74174 30658 74226
rect 31390 74174 31442 74226
rect 32174 74174 32226 74226
rect 36766 74174 36818 74226
rect 37886 74174 37938 74226
rect 38334 74174 38386 74226
rect 38782 74174 38834 74226
rect 4398 74062 4450 74114
rect 4734 74062 4786 74114
rect 4958 74062 5010 74114
rect 6974 74062 7026 74114
rect 7646 74062 7698 74114
rect 7758 74062 7810 74114
rect 7982 74062 8034 74114
rect 8654 74062 8706 74114
rect 8878 74062 8930 74114
rect 9774 74062 9826 74114
rect 9998 74062 10050 74114
rect 10670 74062 10722 74114
rect 11006 74062 11058 74114
rect 11118 74062 11170 74114
rect 11342 74062 11394 74114
rect 12014 74062 12066 74114
rect 13806 74062 13858 74114
rect 17166 74062 17218 74114
rect 22094 74062 22146 74114
rect 23438 74062 23490 74114
rect 30270 74062 30322 74114
rect 32510 74062 32562 74114
rect 32958 74062 33010 74114
rect 33630 74062 33682 74114
rect 34414 74062 34466 74114
rect 35198 74062 35250 74114
rect 35982 74062 36034 74114
rect 3502 73950 3554 74002
rect 3950 73950 4002 74002
rect 7422 73950 7474 74002
rect 8990 73950 9042 74002
rect 10110 73950 10162 74002
rect 12686 73950 12738 74002
rect 12798 73950 12850 74002
rect 12910 73950 12962 74002
rect 20862 73950 20914 74002
rect 21646 73950 21698 74002
rect 22318 73950 22370 74002
rect 22766 73950 22818 74002
rect 24110 73950 24162 74002
rect 28366 73950 28418 74002
rect 30942 73950 30994 74002
rect 37438 73950 37490 74002
rect 6414 73838 6466 73890
rect 20526 73838 20578 73890
rect 20750 73838 20802 73890
rect 21870 73838 21922 73890
rect 22430 73838 22482 73890
rect 33182 73838 33234 73890
rect 36318 73838 36370 73890
rect 39230 73838 39282 73890
rect 39678 73838 39730 73890
rect 40126 73838 40178 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 1934 73502 1986 73554
rect 2382 73502 2434 73554
rect 7646 73502 7698 73554
rect 23998 73502 24050 73554
rect 35534 73502 35586 73554
rect 36430 73502 36482 73554
rect 37326 73502 37378 73554
rect 4174 73390 4226 73442
rect 6750 73390 6802 73442
rect 8990 73390 9042 73442
rect 10222 73390 10274 73442
rect 14814 73390 14866 73442
rect 18510 73390 18562 73442
rect 19182 73390 19234 73442
rect 29150 73390 29202 73442
rect 30494 73390 30546 73442
rect 32398 73390 32450 73442
rect 36878 73390 36930 73442
rect 4510 73278 4562 73330
rect 5182 73278 5234 73330
rect 5406 73278 5458 73330
rect 6190 73278 6242 73330
rect 6414 73278 6466 73330
rect 7198 73278 7250 73330
rect 7870 73278 7922 73330
rect 8878 73278 8930 73330
rect 10670 73278 10722 73330
rect 11342 73278 11394 73330
rect 13022 73278 13074 73330
rect 14030 73278 14082 73330
rect 17726 73278 17778 73330
rect 17950 73278 18002 73330
rect 18174 73278 18226 73330
rect 19406 73278 19458 73330
rect 20190 73278 20242 73330
rect 23662 73278 23714 73330
rect 23998 73278 24050 73330
rect 24334 73278 24386 73330
rect 28590 73278 28642 73330
rect 29374 73278 29426 73330
rect 29710 73278 29762 73330
rect 29822 73278 29874 73330
rect 31502 73278 31554 73330
rect 33966 73278 34018 73330
rect 2830 73166 2882 73218
rect 3278 73166 3330 73218
rect 3726 73166 3778 73218
rect 4286 73166 4338 73218
rect 6638 73166 6690 73218
rect 7758 73166 7810 73218
rect 11790 73166 11842 73218
rect 12798 73166 12850 73218
rect 16942 73166 16994 73218
rect 20862 73166 20914 73218
rect 22990 73166 23042 73218
rect 24894 73166 24946 73218
rect 25678 73166 25730 73218
rect 27806 73166 27858 73218
rect 31726 73166 31778 73218
rect 32846 73166 32898 73218
rect 33742 73166 33794 73218
rect 34638 73166 34690 73218
rect 35086 73166 35138 73218
rect 35982 73166 36034 73218
rect 37774 73166 37826 73218
rect 38222 73166 38274 73218
rect 38670 73166 38722 73218
rect 39118 73166 39170 73218
rect 39566 73166 39618 73218
rect 5070 73054 5122 73106
rect 5518 73054 5570 73106
rect 8542 73054 8594 73106
rect 8654 73054 8706 73106
rect 10222 73054 10274 73106
rect 13358 73054 13410 73106
rect 18398 73054 18450 73106
rect 29150 73054 29202 73106
rect 30270 73054 30322 73106
rect 35534 73054 35586 73106
rect 35982 73054 36034 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 3390 72718 3442 72770
rect 3838 72718 3890 72770
rect 4510 72718 4562 72770
rect 6302 72718 6354 72770
rect 7086 72718 7138 72770
rect 7422 72718 7474 72770
rect 19742 72718 19794 72770
rect 30270 72718 30322 72770
rect 33966 72718 34018 72770
rect 34638 72718 34690 72770
rect 34974 72718 35026 72770
rect 2046 72606 2098 72658
rect 2942 72606 2994 72658
rect 3390 72606 3442 72658
rect 4286 72606 4338 72658
rect 9998 72606 10050 72658
rect 11678 72606 11730 72658
rect 12014 72606 12066 72658
rect 20414 72606 20466 72658
rect 21646 72606 21698 72658
rect 23774 72606 23826 72658
rect 25118 72606 25170 72658
rect 28030 72606 28082 72658
rect 30494 72606 30546 72658
rect 32062 72606 32114 72658
rect 34638 72606 34690 72658
rect 35646 72606 35698 72658
rect 36430 72606 36482 72658
rect 37886 72606 37938 72658
rect 3838 72494 3890 72546
rect 6862 72494 6914 72546
rect 7982 72494 8034 72546
rect 8206 72494 8258 72546
rect 9102 72494 9154 72546
rect 12238 72494 12290 72546
rect 17390 72494 17442 72546
rect 18286 72494 18338 72546
rect 18510 72494 18562 72546
rect 20302 72494 20354 72546
rect 24446 72494 24498 72546
rect 28814 72494 28866 72546
rect 30718 72494 30770 72546
rect 30830 72494 30882 72546
rect 31838 72494 31890 72546
rect 32622 72494 32674 72546
rect 33518 72494 33570 72546
rect 38334 72494 38386 72546
rect 38782 72494 38834 72546
rect 4734 72382 4786 72434
rect 5966 72382 6018 72434
rect 11006 72382 11058 72434
rect 11118 72382 11170 72434
rect 13694 72382 13746 72434
rect 16718 72382 16770 72434
rect 18062 72382 18114 72434
rect 20638 72382 20690 72434
rect 20862 72382 20914 72434
rect 32958 72382 33010 72434
rect 35982 72382 36034 72434
rect 2494 72270 2546 72322
rect 4846 72270 4898 72322
rect 5070 72270 5122 72322
rect 6190 72270 6242 72322
rect 8542 72270 8594 72322
rect 10782 72270 10834 72322
rect 13806 72270 13858 72322
rect 14478 72270 14530 72322
rect 18398 72270 18450 72322
rect 18622 72270 18674 72322
rect 19518 72270 19570 72322
rect 19630 72270 19682 72322
rect 25790 72270 25842 72322
rect 29598 72270 29650 72322
rect 30382 72270 30434 72322
rect 31502 72270 31554 72322
rect 33630 72270 33682 72322
rect 33854 72270 33906 72322
rect 34190 72270 34242 72322
rect 35086 72270 35138 72322
rect 37438 72270 37490 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 1934 71934 1986 71986
rect 2382 71934 2434 71986
rect 5630 71934 5682 71986
rect 9774 71934 9826 71986
rect 18062 71934 18114 71986
rect 18286 71934 18338 71986
rect 27246 71934 27298 71986
rect 32398 71934 32450 71986
rect 34078 71934 34130 71986
rect 36878 71934 36930 71986
rect 37326 71934 37378 71986
rect 5406 71822 5458 71874
rect 5742 71822 5794 71874
rect 6526 71822 6578 71874
rect 8094 71822 8146 71874
rect 29374 71822 29426 71874
rect 33854 71822 33906 71874
rect 35086 71822 35138 71874
rect 35534 71822 35586 71874
rect 3390 71710 3442 71762
rect 3838 71710 3890 71762
rect 5966 71710 6018 71762
rect 7198 71710 7250 71762
rect 10670 71710 10722 71762
rect 10782 71710 10834 71762
rect 10894 71710 10946 71762
rect 16718 71710 16770 71762
rect 18734 71710 18786 71762
rect 19182 71710 19234 71762
rect 24894 71710 24946 71762
rect 25678 71710 25730 71762
rect 25902 71710 25954 71762
rect 26350 71710 26402 71762
rect 27470 71710 27522 71762
rect 27582 71710 27634 71762
rect 27694 71710 27746 71762
rect 28702 71710 28754 71762
rect 29150 71710 29202 71762
rect 30046 71710 30098 71762
rect 30606 71710 30658 71762
rect 31390 71710 31442 71762
rect 32286 71710 32338 71762
rect 32622 71710 32674 71762
rect 32846 71710 32898 71762
rect 34190 71710 34242 71762
rect 37774 71710 37826 71762
rect 2830 71598 2882 71650
rect 4286 71598 4338 71650
rect 4846 71598 4898 71650
rect 8542 71598 8594 71650
rect 13358 71598 13410 71650
rect 18174 71598 18226 71650
rect 24222 71598 24274 71650
rect 25790 71598 25842 71650
rect 28366 71598 28418 71650
rect 34638 71598 34690 71650
rect 35982 71598 36034 71650
rect 36430 71598 36482 71650
rect 38222 71598 38274 71650
rect 10222 71486 10274 71538
rect 26798 71486 26850 71538
rect 26910 71486 26962 71538
rect 36430 71486 36482 71538
rect 36654 71486 36706 71538
rect 37438 71486 37490 71538
rect 38334 71486 38386 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 5630 71150 5682 71202
rect 7310 71150 7362 71202
rect 13918 71150 13970 71202
rect 25230 71150 25282 71202
rect 26126 71150 26178 71202
rect 26238 71150 26290 71202
rect 28590 71150 28642 71202
rect 29598 71150 29650 71202
rect 29710 71150 29762 71202
rect 30158 71150 30210 71202
rect 2158 71038 2210 71090
rect 2606 71038 2658 71090
rect 3502 71038 3554 71090
rect 3950 71038 4002 71090
rect 4622 71038 4674 71090
rect 11902 71038 11954 71090
rect 12798 71038 12850 71090
rect 21646 71038 21698 71090
rect 23774 71038 23826 71090
rect 27134 71038 27186 71090
rect 28702 71038 28754 71090
rect 32062 71038 32114 71090
rect 35198 71038 35250 71090
rect 35534 71038 35586 71090
rect 36430 71038 36482 71090
rect 37438 71038 37490 71090
rect 4398 70926 4450 70978
rect 5966 70926 6018 70978
rect 6302 70926 6354 70978
rect 6414 70926 6466 70978
rect 6526 70926 6578 70978
rect 7422 70926 7474 70978
rect 11006 70926 11058 70978
rect 12686 70926 12738 70978
rect 14142 70926 14194 70978
rect 14366 70926 14418 70978
rect 15262 70926 15314 70978
rect 24558 70926 24610 70978
rect 25566 70926 25618 70978
rect 27582 70926 27634 70978
rect 29934 70926 29986 70978
rect 30382 70926 30434 70978
rect 31502 70926 31554 70978
rect 31838 70926 31890 70978
rect 32958 70926 33010 70978
rect 33406 70926 33458 70978
rect 33742 70926 33794 70978
rect 34638 70926 34690 70978
rect 7310 70814 7362 70866
rect 10334 70814 10386 70866
rect 13694 70814 13746 70866
rect 19182 70814 19234 70866
rect 25118 70814 25170 70866
rect 25454 70814 25506 70866
rect 26462 70814 26514 70866
rect 28030 70814 28082 70866
rect 2942 70702 2994 70754
rect 4958 70702 5010 70754
rect 8094 70702 8146 70754
rect 12462 70702 12514 70754
rect 12910 70702 12962 70754
rect 14814 70702 14866 70754
rect 32622 70702 32674 70754
rect 33630 70702 33682 70754
rect 34190 70702 34242 70754
rect 35982 70702 36034 70754
rect 37886 70702 37938 70754
rect 38334 70702 38386 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 4398 70366 4450 70418
rect 5630 70366 5682 70418
rect 5854 70366 5906 70418
rect 6750 70366 6802 70418
rect 8318 70366 8370 70418
rect 8542 70366 8594 70418
rect 18174 70366 18226 70418
rect 18846 70366 18898 70418
rect 23886 70366 23938 70418
rect 24110 70366 24162 70418
rect 29486 70366 29538 70418
rect 33742 70366 33794 70418
rect 35646 70366 35698 70418
rect 36430 70366 36482 70418
rect 2494 70254 2546 70306
rect 6862 70254 6914 70306
rect 7086 70254 7138 70306
rect 29598 70254 29650 70306
rect 29822 70254 29874 70306
rect 35086 70254 35138 70306
rect 2046 70142 2098 70194
rect 2270 70142 2322 70194
rect 3838 70142 3890 70194
rect 5182 70142 5234 70194
rect 7198 70142 7250 70194
rect 8206 70142 8258 70194
rect 8766 70142 8818 70194
rect 10110 70142 10162 70194
rect 13470 70142 13522 70194
rect 18174 70142 18226 70194
rect 18510 70142 18562 70194
rect 18734 70142 18786 70194
rect 23102 70142 23154 70194
rect 24334 70142 24386 70194
rect 28590 70142 28642 70194
rect 29150 70142 29202 70194
rect 29374 70142 29426 70194
rect 31054 70142 31106 70194
rect 32062 70142 32114 70194
rect 32286 70142 32338 70194
rect 32622 70142 32674 70194
rect 33518 70142 33570 70194
rect 33854 70142 33906 70194
rect 34078 70142 34130 70194
rect 36990 70142 37042 70194
rect 37326 70142 37378 70194
rect 2382 70030 2434 70082
rect 3054 70030 3106 70082
rect 3390 70030 3442 70082
rect 4734 70030 4786 70082
rect 5742 70030 5794 70082
rect 7310 70030 7362 70082
rect 7534 70030 7586 70082
rect 8430 70030 8482 70082
rect 10782 70030 10834 70082
rect 12910 70030 12962 70082
rect 14254 70030 14306 70082
rect 16382 70030 16434 70082
rect 17614 70030 17666 70082
rect 17950 70030 18002 70082
rect 19518 70030 19570 70082
rect 20190 70030 20242 70082
rect 22430 70030 22482 70082
rect 24222 70030 24274 70082
rect 24894 70030 24946 70082
rect 25678 70030 25730 70082
rect 27806 70030 27858 70082
rect 31166 70030 31218 70082
rect 31502 70030 31554 70082
rect 32174 70030 32226 70082
rect 34638 70030 34690 70082
rect 35982 70030 36034 70082
rect 35982 69918 36034 69970
rect 36654 69918 36706 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 5854 69582 5906 69634
rect 6190 69582 6242 69634
rect 6302 69582 6354 69634
rect 28142 69582 28194 69634
rect 31726 69582 31778 69634
rect 32734 69582 32786 69634
rect 33518 69582 33570 69634
rect 1934 69470 1986 69522
rect 3166 69470 3218 69522
rect 4174 69470 4226 69522
rect 4510 69470 4562 69522
rect 4958 69470 5010 69522
rect 7198 69470 7250 69522
rect 13694 69470 13746 69522
rect 17166 69470 17218 69522
rect 19294 69470 19346 69522
rect 22990 69470 23042 69522
rect 25118 69470 25170 69522
rect 34526 69470 34578 69522
rect 34862 69470 34914 69522
rect 35310 69470 35362 69522
rect 35758 69470 35810 69522
rect 3726 69358 3778 69410
rect 5966 69358 6018 69410
rect 7646 69358 7698 69410
rect 7870 69358 7922 69410
rect 8206 69358 8258 69410
rect 9550 69358 9602 69410
rect 10334 69358 10386 69410
rect 12462 69358 12514 69410
rect 13022 69358 13074 69410
rect 16606 69358 16658 69410
rect 19966 69358 20018 69410
rect 22206 69358 22258 69410
rect 26126 69358 26178 69410
rect 26798 69358 26850 69410
rect 27134 69358 27186 69410
rect 28030 69358 28082 69410
rect 28366 69358 28418 69410
rect 28590 69358 28642 69410
rect 28814 69358 28866 69410
rect 30158 69358 30210 69410
rect 32062 69358 32114 69410
rect 33406 69358 33458 69410
rect 34078 69358 34130 69410
rect 9102 69246 9154 69298
rect 11566 69246 11618 69298
rect 11678 69246 11730 69298
rect 15822 69246 15874 69298
rect 20526 69246 20578 69298
rect 20750 69246 20802 69298
rect 2382 69134 2434 69186
rect 2830 69134 2882 69186
rect 10894 69134 10946 69186
rect 11902 69134 11954 69186
rect 12350 69134 12402 69186
rect 12574 69134 12626 69186
rect 20862 69190 20914 69242
rect 30046 69246 30098 69298
rect 30830 69246 30882 69298
rect 21758 69134 21810 69186
rect 25790 69134 25842 69186
rect 26014 69134 26066 69186
rect 26238 69134 26290 69186
rect 27246 69134 27298 69186
rect 27358 69134 27410 69186
rect 29710 69134 29762 69186
rect 29934 69134 29986 69186
rect 30718 69134 30770 69186
rect 31838 69134 31890 69186
rect 32734 69134 32786 69186
rect 32846 69190 32898 69242
rect 36206 69134 36258 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 5070 68798 5122 68850
rect 9886 68798 9938 68850
rect 18510 68798 18562 68850
rect 24894 68798 24946 68850
rect 26014 68798 26066 68850
rect 26126 68798 26178 68850
rect 32958 68798 33010 68850
rect 33966 68798 34018 68850
rect 4398 68686 4450 68738
rect 9774 68686 9826 68738
rect 21198 68686 21250 68738
rect 25678 68686 25730 68738
rect 30046 68686 30098 68738
rect 32846 68686 32898 68738
rect 33518 68686 33570 68738
rect 2046 68574 2098 68626
rect 2382 68574 2434 68626
rect 8878 68574 8930 68626
rect 10446 68574 10498 68626
rect 16718 68574 16770 68626
rect 18174 68574 18226 68626
rect 18398 68574 18450 68626
rect 19182 68574 19234 68626
rect 25902 68574 25954 68626
rect 26238 68574 26290 68626
rect 27246 68574 27298 68626
rect 27470 68574 27522 68626
rect 28254 68574 28306 68626
rect 29038 68574 29090 68626
rect 31614 68574 31666 68626
rect 32286 68574 32338 68626
rect 32622 68574 32674 68626
rect 2942 68462 2994 68514
rect 3390 68462 3442 68514
rect 3838 68462 3890 68514
rect 5182 68462 5234 68514
rect 6078 68462 6130 68514
rect 8206 68462 8258 68514
rect 11790 68462 11842 68514
rect 28702 68462 28754 68514
rect 31390 68462 31442 68514
rect 34414 68462 34466 68514
rect 34862 68462 34914 68514
rect 35310 68462 35362 68514
rect 4286 68350 4338 68402
rect 5294 68350 5346 68402
rect 10670 68350 10722 68402
rect 10894 68350 10946 68402
rect 11006 68350 11058 68402
rect 18510 68350 18562 68402
rect 26910 68350 26962 68402
rect 29934 68350 29986 68402
rect 30942 68350 30994 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 5518 68014 5570 68066
rect 5742 68014 5794 68066
rect 12462 68014 12514 68066
rect 12798 68014 12850 68066
rect 12910 68014 12962 68066
rect 14030 68014 14082 68066
rect 29598 68014 29650 68066
rect 31726 68014 31778 68066
rect 3726 67902 3778 67954
rect 7198 67902 7250 67954
rect 7982 67902 8034 67954
rect 10222 67902 10274 67954
rect 11678 67902 11730 67954
rect 13806 67902 13858 67954
rect 15710 67902 15762 67954
rect 17166 67902 17218 67954
rect 17838 67902 17890 67954
rect 20078 67902 20130 67954
rect 23550 67902 23602 67954
rect 26014 67902 26066 67954
rect 28142 67902 28194 67954
rect 28814 67902 28866 67954
rect 2830 67790 2882 67842
rect 4174 67790 4226 67842
rect 4622 67790 4674 67842
rect 5966 67790 6018 67842
rect 8430 67790 8482 67842
rect 9326 67790 9378 67842
rect 10110 67790 10162 67842
rect 10334 67790 10386 67842
rect 11454 67790 11506 67842
rect 12574 67790 12626 67842
rect 14254 67790 14306 67842
rect 14478 67790 14530 67842
rect 15598 67790 15650 67842
rect 16270 67790 16322 67842
rect 20750 67790 20802 67842
rect 21758 67790 21810 67842
rect 22094 67790 22146 67842
rect 23438 67790 23490 67842
rect 23662 67790 23714 67842
rect 23886 67790 23938 67842
rect 24446 67790 24498 67842
rect 24782 67790 24834 67842
rect 25342 67790 25394 67842
rect 30718 67790 30770 67842
rect 31614 67790 31666 67842
rect 32398 67790 32450 67842
rect 32734 67790 32786 67842
rect 3278 67678 3330 67730
rect 7870 67678 7922 67730
rect 8206 67678 8258 67730
rect 8990 67678 9042 67730
rect 9550 67678 9602 67730
rect 10558 67678 10610 67730
rect 11230 67678 11282 67730
rect 11790 67678 11842 67730
rect 15710 67678 15762 67730
rect 16606 67678 16658 67730
rect 21646 67678 21698 67730
rect 23214 67678 23266 67730
rect 29934 67678 29986 67730
rect 30606 67678 30658 67730
rect 31726 67678 31778 67730
rect 33966 67678 34018 67730
rect 1934 67566 1986 67618
rect 2382 67566 2434 67618
rect 4958 67566 5010 67618
rect 6078 67566 6130 67618
rect 6302 67566 6354 67618
rect 6862 67566 6914 67618
rect 7086 67566 7138 67618
rect 7310 67566 7362 67618
rect 9102 67566 9154 67618
rect 14366 67566 14418 67618
rect 24558 67566 24610 67618
rect 29710 67566 29762 67618
rect 30382 67566 30434 67618
rect 32510 67566 32562 67618
rect 33070 67566 33122 67618
rect 33518 67566 33570 67618
rect 34414 67566 34466 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 3614 67230 3666 67282
rect 6638 67230 6690 67282
rect 8878 67230 8930 67282
rect 17950 67230 18002 67282
rect 31390 67230 31442 67282
rect 31614 67230 31666 67282
rect 31950 67230 32002 67282
rect 3166 67118 3218 67170
rect 4846 67118 4898 67170
rect 5406 67118 5458 67170
rect 4622 67006 4674 67058
rect 1934 66894 1986 66946
rect 2382 66894 2434 66946
rect 2718 66894 2770 66946
rect 4174 66894 4226 66946
rect 3390 66782 3442 66834
rect 7422 67118 7474 67170
rect 10110 67118 10162 67170
rect 14926 67118 14978 67170
rect 20078 67118 20130 67170
rect 22654 67118 22706 67170
rect 24334 67118 24386 67170
rect 26126 67118 26178 67170
rect 26238 67118 26290 67170
rect 26910 67118 26962 67170
rect 27134 67118 27186 67170
rect 28590 67118 28642 67170
rect 29374 67118 29426 67170
rect 32398 67118 32450 67170
rect 32846 67118 32898 67170
rect 6974 67006 7026 67058
rect 7198 67006 7250 67058
rect 7646 67006 7698 67058
rect 8766 67006 8818 67058
rect 10334 67006 10386 67058
rect 10558 67006 10610 67058
rect 11566 67006 11618 67058
rect 15150 67006 15202 67058
rect 15598 67006 15650 67058
rect 16606 67006 16658 67058
rect 18286 67006 18338 67058
rect 18510 67006 18562 67058
rect 19294 67006 19346 67058
rect 23886 67006 23938 67058
rect 25678 67006 25730 67058
rect 26014 67006 26066 67058
rect 26798 67006 26850 67058
rect 27918 67006 27970 67058
rect 29598 67006 29650 67058
rect 30270 67006 30322 67058
rect 30606 67006 30658 67058
rect 31278 67006 31330 67058
rect 4958 66894 5010 66946
rect 5854 66894 5906 66946
rect 6638 66894 6690 66946
rect 8542 66894 8594 66946
rect 10446 66894 10498 66946
rect 12238 66894 12290 66946
rect 14366 66894 14418 66946
rect 15374 66894 15426 66946
rect 16942 66894 16994 66946
rect 17838 66894 17890 66946
rect 22206 66894 22258 66946
rect 23998 66894 24050 66946
rect 24894 66894 24946 66946
rect 27806 66894 27858 66946
rect 29262 66894 29314 66946
rect 6414 66782 6466 66834
rect 7310 66782 7362 66834
rect 16046 66782 16098 66834
rect 16606 66782 16658 66834
rect 18062 66782 18114 66834
rect 27582 66782 27634 66834
rect 32062 66782 32114 66834
rect 32622 66782 32674 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 5966 66446 6018 66498
rect 6414 66446 6466 66498
rect 8094 66446 8146 66498
rect 9326 66446 9378 66498
rect 28814 66446 28866 66498
rect 29934 66446 29986 66498
rect 2158 66334 2210 66386
rect 2606 66334 2658 66386
rect 4062 66334 4114 66386
rect 4622 66334 4674 66386
rect 6302 66334 6354 66386
rect 6750 66334 6802 66386
rect 9214 66334 9266 66386
rect 11902 66334 11954 66386
rect 13694 66334 13746 66386
rect 19294 66334 19346 66386
rect 20078 66334 20130 66386
rect 20862 66334 20914 66386
rect 22878 66334 22930 66386
rect 23438 66334 23490 66386
rect 29598 66334 29650 66386
rect 30606 66334 30658 66386
rect 31502 66334 31554 66386
rect 32062 66334 32114 66386
rect 3166 66222 3218 66274
rect 10558 66222 10610 66274
rect 12686 66222 12738 66274
rect 16494 66222 16546 66274
rect 17166 66222 17218 66274
rect 18510 66222 18562 66274
rect 19966 66222 20018 66274
rect 22206 66222 22258 66274
rect 22766 66222 22818 66274
rect 26238 66222 26290 66274
rect 26910 66222 26962 66274
rect 27134 66222 27186 66274
rect 27582 66222 27634 66274
rect 28254 66222 28306 66274
rect 31278 66222 31330 66274
rect 3390 66110 3442 66162
rect 6862 66110 6914 66162
rect 7422 66110 7474 66162
rect 8318 66110 8370 66162
rect 11566 66110 11618 66162
rect 15822 66110 15874 66162
rect 17390 66110 17442 66162
rect 17502 66110 17554 66162
rect 18622 66110 18674 66162
rect 25566 66110 25618 66162
rect 28142 66110 28194 66162
rect 28366 66110 28418 66162
rect 29710 66110 29762 66162
rect 5070 65998 5122 66050
rect 5742 65998 5794 66050
rect 7534 65998 7586 66050
rect 8206 65998 8258 66050
rect 9102 65998 9154 66050
rect 9998 65998 10050 66050
rect 12798 65998 12850 66050
rect 13022 65998 13074 66050
rect 17950 65998 18002 66050
rect 18846 65998 18898 66050
rect 27022 65998 27074 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 4846 65550 4898 65602
rect 7422 65606 7474 65658
rect 8094 65662 8146 65714
rect 8318 65662 8370 65714
rect 16382 65662 16434 65714
rect 18174 65662 18226 65714
rect 21534 65662 21586 65714
rect 21646 65662 21698 65714
rect 21758 65662 21810 65714
rect 21870 65662 21922 65714
rect 24894 65662 24946 65714
rect 30494 65662 30546 65714
rect 31054 65662 31106 65714
rect 2270 65438 2322 65490
rect 4062 65438 4114 65490
rect 5406 65438 5458 65490
rect 7310 65494 7362 65546
rect 8206 65550 8258 65602
rect 10222 65550 10274 65602
rect 12462 65550 12514 65602
rect 16270 65550 16322 65602
rect 17726 65550 17778 65602
rect 18622 65550 18674 65602
rect 20190 65550 20242 65602
rect 20302 65550 20354 65602
rect 21310 65550 21362 65602
rect 22542 65550 22594 65602
rect 23550 65550 23602 65602
rect 23886 65550 23938 65602
rect 26686 65550 26738 65602
rect 27358 65550 27410 65602
rect 27918 65550 27970 65602
rect 30606 65550 30658 65602
rect 7646 65438 7698 65490
rect 8766 65438 8818 65490
rect 11230 65438 11282 65490
rect 13806 65438 13858 65490
rect 14814 65438 14866 65490
rect 15598 65438 15650 65490
rect 16606 65438 16658 65490
rect 16718 65438 16770 65490
rect 17950 65438 18002 65490
rect 18286 65438 18338 65490
rect 19182 65438 19234 65490
rect 22766 65438 22818 65490
rect 23438 65438 23490 65490
rect 24222 65438 24274 65490
rect 26014 65438 26066 65490
rect 26462 65438 26514 65490
rect 27694 65438 27746 65490
rect 29486 65438 29538 65490
rect 29710 65438 29762 65490
rect 30270 65438 30322 65490
rect 1822 65326 1874 65378
rect 2718 65326 2770 65378
rect 3054 65326 3106 65378
rect 3614 65326 3666 65378
rect 4510 65326 4562 65378
rect 6302 65326 6354 65378
rect 6750 65326 6802 65378
rect 11118 65326 11170 65378
rect 13470 65326 13522 65378
rect 16270 65326 16322 65378
rect 28814 65326 28866 65378
rect 4510 65214 4562 65266
rect 5182 65214 5234 65266
rect 5518 65214 5570 65266
rect 6526 65214 6578 65266
rect 7086 65214 7138 65266
rect 10110 65214 10162 65266
rect 10446 65214 10498 65266
rect 18174 65214 18226 65266
rect 19742 65214 19794 65266
rect 19966 65214 20018 65266
rect 20526 65214 20578 65266
rect 24446 65214 24498 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 2046 64878 2098 64930
rect 2606 64878 2658 64930
rect 3614 64878 3666 64930
rect 1934 64766 1986 64818
rect 2382 64766 2434 64818
rect 3166 64654 3218 64706
rect 11902 64878 11954 64930
rect 14254 64878 14306 64930
rect 15374 64878 15426 64930
rect 16046 64878 16098 64930
rect 27022 64878 27074 64930
rect 4958 64766 5010 64818
rect 6078 64766 6130 64818
rect 14030 64766 14082 64818
rect 17726 64766 17778 64818
rect 20526 64766 20578 64818
rect 22094 64766 22146 64818
rect 23102 64766 23154 64818
rect 23998 64766 24050 64818
rect 27470 64766 27522 64818
rect 28254 64766 28306 64818
rect 29822 64766 29874 64818
rect 30270 64766 30322 64818
rect 3614 64654 3666 64706
rect 4846 64654 4898 64706
rect 7534 64654 7586 64706
rect 9438 64654 9490 64706
rect 14366 64654 14418 64706
rect 15486 64654 15538 64706
rect 15710 64654 15762 64706
rect 15934 64654 15986 64706
rect 16830 64654 16882 64706
rect 17166 64654 17218 64706
rect 18958 64654 19010 64706
rect 19854 64654 19906 64706
rect 20190 64654 20242 64706
rect 23774 64654 23826 64706
rect 23886 64654 23938 64706
rect 24110 64654 24162 64706
rect 24334 64654 24386 64706
rect 25118 64654 25170 64706
rect 25342 64654 25394 64706
rect 26350 64654 26402 64706
rect 26686 64654 26738 64706
rect 28030 64654 28082 64706
rect 2830 64542 2882 64594
rect 4510 64542 4562 64594
rect 6526 64542 6578 64594
rect 9662 64542 9714 64594
rect 9774 64542 9826 64594
rect 9998 64542 10050 64594
rect 12126 64542 12178 64594
rect 12574 64542 12626 64594
rect 18398 64542 18450 64594
rect 25678 64542 25730 64594
rect 26910 64542 26962 64594
rect 4062 64430 4114 64482
rect 7870 64430 7922 64482
rect 8990 64430 9042 64482
rect 9550 64430 9602 64482
rect 10894 64430 10946 64482
rect 11566 64430 11618 64482
rect 18286 64430 18338 64482
rect 18510 64430 18562 64482
rect 20862 64430 20914 64482
rect 21982 64430 22034 64482
rect 22206 64430 22258 64482
rect 22430 64430 22482 64482
rect 25566 64430 25618 64482
rect 25790 64430 25842 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 1934 64094 1986 64146
rect 2718 64094 2770 64146
rect 4622 64094 4674 64146
rect 5518 64094 5570 64146
rect 5854 64094 5906 64146
rect 7198 64094 7250 64146
rect 8206 64094 8258 64146
rect 11454 64094 11506 64146
rect 12126 64094 12178 64146
rect 15038 64094 15090 64146
rect 15150 64094 15202 64146
rect 15262 64094 15314 64146
rect 16382 64094 16434 64146
rect 16494 64094 16546 64146
rect 16606 64094 16658 64146
rect 18174 64094 18226 64146
rect 19182 64094 19234 64146
rect 20302 64094 20354 64146
rect 20526 64094 20578 64146
rect 22766 64094 22818 64146
rect 24110 64094 24162 64146
rect 24894 64094 24946 64146
rect 26798 64094 26850 64146
rect 27806 64094 27858 64146
rect 28590 64094 28642 64146
rect 28926 64094 28978 64146
rect 12350 63982 12402 64034
rect 19070 63982 19122 64034
rect 19630 63982 19682 64034
rect 20190 63982 20242 64034
rect 23326 63982 23378 64034
rect 25790 63982 25842 64034
rect 25902 63982 25954 64034
rect 2382 63870 2434 63922
rect 3726 63870 3778 63922
rect 6302 63870 6354 63922
rect 6862 63870 6914 63922
rect 8766 63870 8818 63922
rect 9998 63870 10050 63922
rect 12014 63870 12066 63922
rect 12574 63870 12626 63922
rect 13582 63870 13634 63922
rect 15486 63870 15538 63922
rect 16942 63870 16994 63922
rect 18062 63870 18114 63922
rect 18398 63870 18450 63922
rect 19294 63870 19346 63922
rect 21534 63870 21586 63922
rect 22206 63870 22258 63922
rect 25566 63870 25618 63922
rect 26686 63870 26738 63922
rect 26910 63870 26962 63922
rect 27358 63870 27410 63922
rect 3166 63758 3218 63810
rect 4062 63758 4114 63810
rect 4958 63758 5010 63810
rect 7646 63758 7698 63810
rect 10334 63758 10386 63810
rect 13918 63758 13970 63810
rect 17726 63758 17778 63810
rect 18286 63758 18338 63810
rect 21310 63758 21362 63810
rect 1710 63646 1762 63698
rect 2830 63646 2882 63698
rect 4062 63646 4114 63698
rect 6862 63646 6914 63698
rect 8542 63646 8594 63698
rect 13694 63646 13746 63698
rect 15710 63646 15762 63698
rect 23886 63646 23938 63698
rect 24222 63646 24274 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 2494 63310 2546 63362
rect 3278 63310 3330 63362
rect 4510 63310 4562 63362
rect 6526 63310 6578 63362
rect 8654 63310 8706 63362
rect 10334 63310 10386 63362
rect 15934 63310 15986 63362
rect 19742 63310 19794 63362
rect 22878 63310 22930 63362
rect 24334 63310 24386 63362
rect 25118 63310 25170 63362
rect 1934 63198 1986 63250
rect 2718 63198 2770 63250
rect 3166 63198 3218 63250
rect 3614 63198 3666 63250
rect 4174 63198 4226 63250
rect 4622 63198 4674 63250
rect 6526 63198 6578 63250
rect 6862 63198 6914 63250
rect 8206 63198 8258 63250
rect 9998 63198 10050 63250
rect 10558 63198 10610 63250
rect 12014 63198 12066 63250
rect 12910 63198 12962 63250
rect 15262 63198 15314 63250
rect 16046 63198 16098 63250
rect 17614 63198 17666 63250
rect 18398 63198 18450 63250
rect 20414 63198 20466 63250
rect 22990 63198 23042 63250
rect 23662 63198 23714 63250
rect 25902 63198 25954 63250
rect 27246 63198 27298 63250
rect 27694 63198 27746 63250
rect 28814 63198 28866 63250
rect 2382 63086 2434 63138
rect 7870 63086 7922 63138
rect 8654 63086 8706 63138
rect 9214 63086 9266 63138
rect 11342 63086 11394 63138
rect 12238 63086 12290 63138
rect 13806 63086 13858 63138
rect 14366 63086 14418 63138
rect 16718 63086 16770 63138
rect 17502 63086 17554 63138
rect 18622 63086 18674 63138
rect 21758 63086 21810 63138
rect 21870 63086 21922 63138
rect 22318 63086 22370 63138
rect 24222 63086 24274 63138
rect 25230 63086 25282 63138
rect 29934 63086 29986 63138
rect 13694 62974 13746 63026
rect 17614 62974 17666 63026
rect 19630 62974 19682 63026
rect 19742 62974 19794 63026
rect 25118 62974 25170 63026
rect 28478 62974 28530 63026
rect 29598 62974 29650 63026
rect 4958 62862 5010 62914
rect 6078 62862 6130 62914
rect 7310 62862 7362 62914
rect 9326 62862 9378 62914
rect 9550 62862 9602 62914
rect 20862 62862 20914 62914
rect 21982 62862 22034 62914
rect 22094 62862 22146 62914
rect 24334 62862 24386 62914
rect 26350 62862 26402 62914
rect 26798 62862 26850 62914
rect 29710 62862 29762 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 1934 62526 1986 62578
rect 2382 62526 2434 62578
rect 2718 62526 2770 62578
rect 3278 62526 3330 62578
rect 3614 62526 3666 62578
rect 4510 62526 4562 62578
rect 5518 62526 5570 62578
rect 5966 62526 6018 62578
rect 6414 62526 6466 62578
rect 7198 62526 7250 62578
rect 7758 62526 7810 62578
rect 8542 62526 8594 62578
rect 8990 62526 9042 62578
rect 10782 62526 10834 62578
rect 12238 62526 12290 62578
rect 13358 62526 13410 62578
rect 13470 62526 13522 62578
rect 13694 62526 13746 62578
rect 15038 62526 15090 62578
rect 15262 62526 15314 62578
rect 15822 62526 15874 62578
rect 16494 62526 16546 62578
rect 16718 62526 16770 62578
rect 19742 62526 19794 62578
rect 20190 62526 20242 62578
rect 20638 62526 20690 62578
rect 21086 62526 21138 62578
rect 21534 62526 21586 62578
rect 22766 62526 22818 62578
rect 23326 62526 23378 62578
rect 23774 62526 23826 62578
rect 24334 62526 24386 62578
rect 24670 62526 24722 62578
rect 25566 62526 25618 62578
rect 26126 62526 26178 62578
rect 26686 62526 26738 62578
rect 27582 62526 27634 62578
rect 28254 62526 28306 62578
rect 28814 62526 28866 62578
rect 11678 62414 11730 62466
rect 15934 62414 15986 62466
rect 22094 62414 22146 62466
rect 22206 62414 22258 62466
rect 28366 62414 28418 62466
rect 4846 62302 4898 62354
rect 4958 62302 5010 62354
rect 4174 62190 4226 62242
rect 8094 62302 8146 62354
rect 10558 62302 10610 62354
rect 11230 62302 11282 62354
rect 11902 62302 11954 62354
rect 13582 62302 13634 62354
rect 13918 62302 13970 62354
rect 14926 62302 14978 62354
rect 16830 62302 16882 62354
rect 28030 62302 28082 62354
rect 6750 62190 6802 62242
rect 9998 62190 10050 62242
rect 10670 62190 10722 62242
rect 12686 62190 12738 62242
rect 14366 62190 14418 62242
rect 17950 62190 18002 62242
rect 19294 62190 19346 62242
rect 8430 62078 8482 62130
rect 12462 62078 12514 62130
rect 12686 62078 12738 62130
rect 15710 62078 15762 62130
rect 18174 62078 18226 62130
rect 18510 62078 18562 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 3390 61742 3442 61794
rect 4062 61742 4114 61794
rect 6302 61742 6354 61794
rect 6750 61742 6802 61794
rect 7422 61742 7474 61794
rect 12574 61742 12626 61794
rect 12910 61742 12962 61794
rect 15710 61742 15762 61794
rect 16158 61742 16210 61794
rect 17278 61742 17330 61794
rect 17502 61742 17554 61794
rect 17950 61742 18002 61794
rect 21870 61742 21922 61794
rect 22430 61742 22482 61794
rect 2382 61630 2434 61682
rect 2718 61630 2770 61682
rect 3166 61630 3218 61682
rect 4510 61630 4562 61682
rect 4958 61630 5010 61682
rect 5854 61630 5906 61682
rect 6302 61630 6354 61682
rect 7198 61630 7250 61682
rect 7758 61630 7810 61682
rect 8878 61630 8930 61682
rect 9326 61630 9378 61682
rect 9886 61630 9938 61682
rect 10782 61630 10834 61682
rect 10894 61630 10946 61682
rect 11566 61630 11618 61682
rect 13806 61630 13858 61682
rect 17166 61630 17218 61682
rect 20750 61630 20802 61682
rect 21758 61630 21810 61682
rect 22206 61630 22258 61682
rect 23550 61630 23602 61682
rect 24222 61630 24274 61682
rect 25006 61630 25058 61682
rect 25342 61630 25394 61682
rect 25902 61630 25954 61682
rect 4062 61518 4114 61570
rect 6750 61518 6802 61570
rect 10222 61518 10274 61570
rect 11118 61518 11170 61570
rect 12574 61518 12626 61570
rect 14366 61518 14418 61570
rect 15150 61518 15202 61570
rect 15822 61518 15874 61570
rect 16046 61518 16098 61570
rect 19742 61518 19794 61570
rect 14702 61406 14754 61458
rect 16718 61406 16770 61458
rect 1934 61294 1986 61346
rect 3614 61294 3666 61346
rect 8430 61294 8482 61346
rect 12014 61294 12066 61346
rect 13694 61294 13746 61346
rect 13918 61294 13970 61346
rect 17614 61294 17666 61346
rect 18062 61294 18114 61346
rect 18734 61294 18786 61346
rect 19182 61294 19234 61346
rect 20302 61294 20354 61346
rect 22654 61294 22706 61346
rect 23102 61294 23154 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 1934 60958 1986 61010
rect 2382 60958 2434 61010
rect 2830 60958 2882 61010
rect 3166 60958 3218 61010
rect 4174 60958 4226 61010
rect 4958 60958 5010 61010
rect 5854 60958 5906 61010
rect 6862 60958 6914 61010
rect 8654 60958 8706 61010
rect 10110 60958 10162 61010
rect 10222 60958 10274 61010
rect 10782 60958 10834 61010
rect 13470 60958 13522 61010
rect 13694 60958 13746 61010
rect 14478 60958 14530 61010
rect 15038 60958 15090 61010
rect 15374 60958 15426 61010
rect 17054 60958 17106 61010
rect 18286 60958 18338 61010
rect 19742 60958 19794 61010
rect 20638 60958 20690 61010
rect 21870 60958 21922 61010
rect 22318 60958 22370 61010
rect 22654 60958 22706 61010
rect 23550 60958 23602 61010
rect 24110 60958 24162 61010
rect 29822 60958 29874 61010
rect 30382 60958 30434 61010
rect 30942 60958 30994 61010
rect 7758 60846 7810 60898
rect 13358 60846 13410 60898
rect 14030 60846 14082 60898
rect 15822 60846 15874 60898
rect 17614 60846 17666 60898
rect 30270 60846 30322 60898
rect 5518 60734 5570 60786
rect 6302 60734 6354 60786
rect 19182 60734 19234 60786
rect 3726 60622 3778 60674
rect 4510 60622 4562 60674
rect 7198 60622 7250 60674
rect 8094 60622 8146 60674
rect 8990 60622 9042 60674
rect 11454 60622 11506 60674
rect 11902 60622 11954 60674
rect 12350 60622 12402 60674
rect 12798 60622 12850 60674
rect 16270 60622 16322 60674
rect 18734 60622 18786 60674
rect 20190 60622 20242 60674
rect 21310 60622 21362 60674
rect 23214 60622 23266 60674
rect 9998 60510 10050 60562
rect 18734 60510 18786 60562
rect 19406 60510 19458 60562
rect 30382 60510 30434 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 3502 60174 3554 60226
rect 4846 60174 4898 60226
rect 2158 60062 2210 60114
rect 2606 60062 2658 60114
rect 3054 60062 3106 60114
rect 3390 60062 3442 60114
rect 3950 60062 4002 60114
rect 4846 60062 4898 60114
rect 7758 60062 7810 60114
rect 8206 60062 8258 60114
rect 8654 60062 8706 60114
rect 8990 60062 9042 60114
rect 9438 60062 9490 60114
rect 10670 60062 10722 60114
rect 11230 60062 11282 60114
rect 12686 60062 12738 60114
rect 13582 60062 13634 60114
rect 14254 60062 14306 60114
rect 14702 60062 14754 60114
rect 15822 60062 15874 60114
rect 16382 60062 16434 60114
rect 16830 60062 16882 60114
rect 17614 60062 17666 60114
rect 19518 60062 19570 60114
rect 20414 60062 20466 60114
rect 20862 60062 20914 60114
rect 21982 60062 22034 60114
rect 23214 60062 23266 60114
rect 23662 60062 23714 60114
rect 6302 59950 6354 60002
rect 11678 59950 11730 60002
rect 18286 59950 18338 60002
rect 9998 59838 10050 59890
rect 15374 59838 15426 59890
rect 19070 59838 19122 59890
rect 4398 59726 4450 59778
rect 5854 59726 5906 59778
rect 6638 59726 6690 59778
rect 7086 59726 7138 59778
rect 17278 59726 17330 59778
rect 19854 59726 19906 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 3950 59390 4002 59442
rect 4734 59390 4786 59442
rect 5294 59390 5346 59442
rect 6302 59390 6354 59442
rect 6862 59390 6914 59442
rect 7310 59390 7362 59442
rect 8654 59390 8706 59442
rect 9102 59390 9154 59442
rect 9774 59390 9826 59442
rect 11230 59390 11282 59442
rect 11678 59390 11730 59442
rect 12462 59390 12514 59442
rect 13022 59390 13074 59442
rect 14926 59390 14978 59442
rect 15486 59390 15538 59442
rect 15934 59390 15986 59442
rect 16494 59390 16546 59442
rect 16942 59390 16994 59442
rect 17726 59390 17778 59442
rect 18510 59390 18562 59442
rect 13582 59278 13634 59330
rect 3390 59054 3442 59106
rect 4398 59054 4450 59106
rect 5966 59054 6018 59106
rect 7646 59054 7698 59106
rect 8094 59054 8146 59106
rect 10446 59054 10498 59106
rect 10782 59054 10834 59106
rect 14030 59054 14082 59106
rect 18174 59054 18226 59106
rect 18958 59054 19010 59106
rect 6078 58942 6130 58994
rect 6638 58942 6690 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 15598 58606 15650 58658
rect 16270 58606 16322 58658
rect 19518 58606 19570 58658
rect 4062 58494 4114 58546
rect 5854 58494 5906 58546
rect 6302 58494 6354 58546
rect 9326 58494 9378 58546
rect 9774 58494 9826 58546
rect 10222 58494 10274 58546
rect 11230 58494 11282 58546
rect 11678 58494 11730 58546
rect 12126 58494 12178 58546
rect 12574 58494 12626 58546
rect 13022 58494 13074 58546
rect 13694 58494 13746 58546
rect 15038 58494 15090 58546
rect 15374 58494 15426 58546
rect 15934 58494 15986 58546
rect 16270 58494 16322 58546
rect 17166 58494 17218 58546
rect 17726 58494 17778 58546
rect 18174 58494 18226 58546
rect 19630 58494 19682 58546
rect 20078 58494 20130 58546
rect 10670 58382 10722 58434
rect 6750 58158 6802 58210
rect 7198 58158 7250 58210
rect 7646 58158 7698 58210
rect 8094 58158 8146 58210
rect 8766 58158 8818 58210
rect 14030 58158 14082 58210
rect 14478 58158 14530 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 7870 57822 7922 57874
rect 8318 57822 8370 57874
rect 8990 57822 9042 57874
rect 9774 57822 9826 57874
rect 10446 57822 10498 57874
rect 11118 57822 11170 57874
rect 11566 57822 11618 57874
rect 12014 57822 12066 57874
rect 12462 57822 12514 57874
rect 13022 57822 13074 57874
rect 15150 57822 15202 57874
rect 13806 57710 13858 57762
rect 14254 57598 14306 57650
rect 7310 57486 7362 57538
rect 13358 57486 13410 57538
rect 14702 57486 14754 57538
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 9326 56926 9378 56978
rect 9774 56926 9826 56978
rect 10222 56926 10274 56978
rect 14142 56926 14194 56978
rect 13582 56814 13634 56866
rect 12574 56590 12626 56642
rect 12910 56590 12962 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 28814 55246 28866 55298
rect 29598 55246 29650 55298
rect 29934 55022 29986 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 17614 36654 17666 36706
rect 16942 36542 16994 36594
rect 17502 36430 17554 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 12462 6078 12514 6130
rect 14366 6078 14418 6130
rect 14814 6078 14866 6130
rect 51214 6078 51266 6130
rect 19630 5966 19682 6018
rect 11006 5854 11058 5906
rect 18622 5854 18674 5906
rect 52222 5854 52274 5906
rect 12126 5742 12178 5794
rect 15374 5742 15426 5794
rect 18174 5742 18226 5794
rect 34302 5742 34354 5794
rect 51774 5742 51826 5794
rect 11230 5630 11282 5682
rect 11566 5630 11618 5682
rect 18846 5630 18898 5682
rect 19182 5630 19234 5682
rect 52446 5630 52498 5682
rect 52782 5630 52834 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 22766 5182 22818 5234
rect 23214 5182 23266 5234
rect 32622 5182 32674 5234
rect 33070 5182 33122 5234
rect 34302 5182 34354 5234
rect 34750 5182 34802 5234
rect 40014 5182 40066 5234
rect 40462 5182 40514 5234
rect 46846 5182 46898 5234
rect 47742 5182 47794 5234
rect 53342 5182 53394 5234
rect 11454 5070 11506 5122
rect 22206 5070 22258 5122
rect 23438 5070 23490 5122
rect 32062 5070 32114 5122
rect 33294 5070 33346 5122
rect 34974 5070 35026 5122
rect 39454 5070 39506 5122
rect 40686 5070 40738 5122
rect 47182 5070 47234 5122
rect 47966 5070 48018 5122
rect 52334 5070 52386 5122
rect 23774 4958 23826 5010
rect 24334 4958 24386 5010
rect 11678 4846 11730 4898
rect 24670 4846 24722 4898
rect 33630 4846 33682 4898
rect 35310 4846 35362 4898
rect 41022 4846 41074 4898
rect 48302 4846 48354 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 12350 4510 12402 4562
rect 14590 4510 14642 4562
rect 26798 4510 26850 4562
rect 27246 4510 27298 4562
rect 50766 4510 50818 4562
rect 51214 4510 51266 4562
rect 7310 4398 7362 4450
rect 12798 4398 12850 4450
rect 16606 4398 16658 4450
rect 19630 4398 19682 4450
rect 19966 4398 20018 4450
rect 29598 4398 29650 4450
rect 34302 4398 34354 4450
rect 34638 4398 34690 4450
rect 38334 4398 38386 4450
rect 38670 4398 38722 4450
rect 43486 4398 43538 4450
rect 43822 4398 43874 4450
rect 49534 4398 49586 4450
rect 49870 4398 49922 4450
rect 54350 4398 54402 4450
rect 54910 4398 54962 4450
rect 55246 4398 55298 4450
rect 58270 4398 58322 4450
rect 66222 4398 66274 4450
rect 7646 4286 7698 4338
rect 11342 4286 11394 4338
rect 11678 4286 11730 4338
rect 11902 4286 11954 4338
rect 15150 4286 15202 4338
rect 15374 4286 15426 4338
rect 15710 4286 15762 4338
rect 16270 4286 16322 4338
rect 27806 4286 27858 4338
rect 28030 4286 28082 4338
rect 28366 4286 28418 4338
rect 29262 4286 29314 4338
rect 51774 4286 51826 4338
rect 51998 4286 52050 4338
rect 52894 4286 52946 4338
rect 53118 4286 53170 4338
rect 53454 4286 53506 4338
rect 54014 4286 54066 4338
rect 57934 4286 57986 4338
rect 65886 4286 65938 4338
rect 74398 4286 74450 4338
rect 75182 4286 75234 4338
rect 52334 4174 52386 4226
rect 65326 4174 65378 4226
rect 76078 4174 76130 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 53006 3726 53058 3778
rect 7870 3614 7922 3666
rect 12238 3614 12290 3666
rect 16046 3614 16098 3666
rect 18174 3614 18226 3666
rect 22094 3614 22146 3666
rect 26686 3614 26738 3666
rect 31390 3614 31442 3666
rect 35758 3614 35810 3666
rect 41694 3614 41746 3666
rect 45614 3614 45666 3666
rect 52110 3614 52162 3666
rect 54910 3614 54962 3666
rect 59278 3614 59330 3666
rect 65214 3614 65266 3666
rect 69134 3614 69186 3666
rect 73726 3614 73778 3666
rect 3502 3502 3554 3554
rect 4286 3502 4338 3554
rect 7310 3502 7362 3554
rect 11566 3502 11618 3554
rect 17502 3502 17554 3554
rect 21422 3502 21474 3554
rect 26014 3502 26066 3554
rect 30718 3502 30770 3554
rect 35086 3502 35138 3554
rect 41022 3502 41074 3554
rect 44942 3502 44994 3554
rect 50542 3502 50594 3554
rect 51662 3502 51714 3554
rect 52782 3502 52834 3554
rect 53342 3502 53394 3554
rect 54350 3502 54402 3554
rect 58606 3502 58658 3554
rect 64542 3502 64594 3554
rect 68462 3502 68514 3554
rect 72606 3502 72658 3554
rect 73278 3502 73330 3554
rect 2606 3390 2658 3442
rect 49646 3390 49698 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2268 79212 2660 79268
rect 2044 78820 2100 78830
rect 2044 76690 2100 78764
rect 2044 76638 2046 76690
rect 2098 76638 2100 76690
rect 2044 76626 2100 76638
rect 2156 77364 2212 77374
rect 2044 76468 2100 76478
rect 2044 75908 2100 76412
rect 2044 75776 2100 75852
rect 2044 75460 2100 75470
rect 1932 74788 1988 74798
rect 1820 74786 1988 74788
rect 1820 74734 1934 74786
rect 1986 74734 1988 74786
rect 1820 74732 1988 74734
rect 1596 74676 1652 74686
rect 1596 60116 1652 74620
rect 1708 70644 1764 70654
rect 1708 63698 1764 70588
rect 1820 69524 1876 74732
rect 1932 74722 1988 74732
rect 2044 74004 2100 75404
rect 2156 74226 2212 77308
rect 2156 74174 2158 74226
rect 2210 74174 2212 74226
rect 2156 74162 2212 74174
rect 2044 73948 2212 74004
rect 1932 73556 1988 73566
rect 1932 73462 1988 73500
rect 2044 72660 2100 72670
rect 2044 72566 2100 72604
rect 1932 72212 1988 72222
rect 1932 71986 1988 72156
rect 1932 71934 1934 71986
rect 1986 71934 1988 71986
rect 1932 71922 1988 71934
rect 2156 71316 2212 73948
rect 2044 71260 2212 71316
rect 2044 70194 2100 71260
rect 2156 71092 2212 71102
rect 2268 71092 2324 79212
rect 2380 79044 2436 79054
rect 2604 79044 2660 79212
rect 2800 79200 2912 80000
rect 3052 79940 3108 79950
rect 2828 79044 2884 79200
rect 2604 78988 2884 79044
rect 2380 75122 2436 78988
rect 2940 78596 2996 78606
rect 2716 77924 2772 77934
rect 2492 77812 2548 77822
rect 2492 76690 2548 77756
rect 2492 76638 2494 76690
rect 2546 76638 2548 76690
rect 2492 76626 2548 76638
rect 2380 75070 2382 75122
rect 2434 75070 2436 75122
rect 2380 75058 2436 75070
rect 2604 75572 2660 75582
rect 2380 74340 2436 74350
rect 2380 73554 2436 74284
rect 2604 74226 2660 75516
rect 2604 74174 2606 74226
rect 2658 74174 2660 74226
rect 2604 74162 2660 74174
rect 2716 74004 2772 77868
rect 2940 76690 2996 78540
rect 2940 76638 2942 76690
rect 2994 76638 2996 76690
rect 2940 76626 2996 76638
rect 2828 75460 2884 75470
rect 2828 75366 2884 75404
rect 2828 74676 2884 74686
rect 2828 74582 2884 74620
rect 2940 74338 2996 74350
rect 2940 74286 2942 74338
rect 2994 74286 2996 74338
rect 2380 73502 2382 73554
rect 2434 73502 2436 73554
rect 2380 73490 2436 73502
rect 2604 73948 2772 74004
rect 2828 74228 2884 74238
rect 2492 72322 2548 72334
rect 2492 72270 2494 72322
rect 2546 72270 2548 72322
rect 2380 71988 2436 71998
rect 2380 71894 2436 71932
rect 2156 71090 2324 71092
rect 2156 71038 2158 71090
rect 2210 71038 2324 71090
rect 2156 71036 2324 71038
rect 2156 71026 2212 71036
rect 2268 70868 2324 71036
rect 2268 70802 2324 70812
rect 2380 70644 2436 70654
rect 2044 70142 2046 70194
rect 2098 70142 2100 70194
rect 1932 69524 1988 69534
rect 1820 69468 1932 69524
rect 1932 69392 1988 69468
rect 2044 68852 2100 70142
rect 2268 70420 2324 70430
rect 2268 70194 2324 70364
rect 2380 70308 2436 70588
rect 2492 70532 2548 72270
rect 2604 71090 2660 73948
rect 2828 73444 2884 74172
rect 2940 73948 2996 74286
rect 3052 74226 3108 79884
rect 4956 79492 5012 79502
rect 4508 79156 4564 79166
rect 4172 79044 4228 79054
rect 3836 78708 3892 78718
rect 3388 78372 3444 78382
rect 3276 76804 3332 76814
rect 3164 74900 3220 74910
rect 3276 74900 3332 76748
rect 3388 76020 3444 78316
rect 3500 76580 3556 76590
rect 3500 76486 3556 76524
rect 3612 76466 3668 76478
rect 3612 76414 3614 76466
rect 3666 76414 3668 76466
rect 3388 75954 3444 75964
rect 3500 76356 3556 76366
rect 3500 75796 3556 76300
rect 3612 76244 3668 76414
rect 3612 76178 3668 76188
rect 3724 76242 3780 76254
rect 3724 76190 3726 76242
rect 3778 76190 3780 76242
rect 3164 74898 3332 74900
rect 3164 74846 3166 74898
rect 3218 74846 3332 74898
rect 3164 74844 3332 74846
rect 3164 74834 3220 74844
rect 3052 74174 3054 74226
rect 3106 74174 3108 74226
rect 3052 74162 3108 74174
rect 3164 74674 3220 74686
rect 3164 74622 3166 74674
rect 3218 74622 3220 74674
rect 2940 73892 3108 73948
rect 2828 73388 2996 73444
rect 2828 73220 2884 73230
rect 2828 73126 2884 73164
rect 2940 72658 2996 73388
rect 2940 72606 2942 72658
rect 2994 72606 2996 72658
rect 2940 72594 2996 72606
rect 2828 71652 2884 71662
rect 2828 71558 2884 71596
rect 2604 71038 2606 71090
rect 2658 71038 2660 71090
rect 2604 71026 2660 71038
rect 2940 70756 2996 70766
rect 2716 70754 2996 70756
rect 2716 70702 2942 70754
rect 2994 70702 2996 70754
rect 2716 70700 2996 70702
rect 2492 70476 2660 70532
rect 2492 70308 2548 70318
rect 2380 70306 2548 70308
rect 2380 70254 2494 70306
rect 2546 70254 2548 70306
rect 2380 70252 2548 70254
rect 2492 70242 2548 70252
rect 2268 70142 2270 70194
rect 2322 70142 2324 70194
rect 2268 70130 2324 70142
rect 2380 70084 2436 70094
rect 2380 69990 2436 70028
rect 1932 68796 2100 68852
rect 2156 69300 2212 69310
rect 1932 68068 1988 68796
rect 2044 68628 2100 68638
rect 2044 68534 2100 68572
rect 1932 68002 1988 68012
rect 1932 67620 1988 67630
rect 1932 67526 1988 67564
rect 2044 67508 2100 67518
rect 1932 66946 1988 66958
rect 1932 66894 1934 66946
rect 1986 66894 1988 66946
rect 1932 65940 1988 66894
rect 1932 65874 1988 65884
rect 1932 65604 1988 65614
rect 1820 65378 1876 65390
rect 1820 65326 1822 65378
rect 1874 65326 1876 65378
rect 1820 64036 1876 65326
rect 1932 64818 1988 65548
rect 1932 64766 1934 64818
rect 1986 64766 1988 64818
rect 1932 64754 1988 64766
rect 2044 64930 2100 67452
rect 2044 64878 2046 64930
rect 2098 64878 2100 64930
rect 1932 64148 1988 64158
rect 2044 64148 2100 64878
rect 1932 64146 2100 64148
rect 1932 64094 1934 64146
rect 1986 64094 2100 64146
rect 1932 64092 2100 64094
rect 2156 66386 2212 69244
rect 2380 69186 2436 69198
rect 2380 69134 2382 69186
rect 2434 69134 2436 69186
rect 2380 68852 2436 69134
rect 2380 68786 2436 68796
rect 2492 69188 2548 69198
rect 2380 68628 2436 68638
rect 2492 68628 2548 69132
rect 2380 68626 2548 68628
rect 2380 68574 2382 68626
rect 2434 68574 2548 68626
rect 2380 68572 2548 68574
rect 2380 68562 2436 68572
rect 2380 67618 2436 67630
rect 2380 67566 2382 67618
rect 2434 67566 2436 67618
rect 2380 67396 2436 67566
rect 2380 67330 2436 67340
rect 2604 67172 2660 70476
rect 2716 67172 2772 70700
rect 2940 70690 2996 70700
rect 3052 70308 3108 73892
rect 2940 70252 3108 70308
rect 2828 69186 2884 69198
rect 2828 69134 2830 69186
rect 2882 69134 2884 69186
rect 2828 69076 2884 69134
rect 2828 69010 2884 69020
rect 2940 68740 2996 70252
rect 3052 70082 3108 70094
rect 3052 70030 3054 70082
rect 3106 70030 3108 70082
rect 3052 69972 3108 70030
rect 3052 69906 3108 69916
rect 3164 69860 3220 74622
rect 3276 74338 3332 74844
rect 3276 74286 3278 74338
rect 3330 74286 3332 74338
rect 3276 74274 3332 74286
rect 3388 75740 3556 75796
rect 3612 76020 3668 76030
rect 3612 75794 3668 75964
rect 3612 75742 3614 75794
rect 3666 75742 3668 75794
rect 3388 73556 3444 75740
rect 3612 75730 3668 75742
rect 3724 75796 3780 76190
rect 3724 75730 3780 75740
rect 3724 75572 3780 75582
rect 3724 75236 3780 75516
rect 3836 75460 3892 78652
rect 4060 77476 4116 77486
rect 3948 76692 4004 76702
rect 3948 75572 4004 76636
rect 4060 75738 4116 77420
rect 4060 75686 4062 75738
rect 4114 75686 4116 75738
rect 4060 75674 4116 75686
rect 4172 75572 4228 78988
rect 4396 76468 4452 76478
rect 4396 76374 4452 76412
rect 4508 76356 4564 79100
rect 4844 78484 4900 78494
rect 4620 77588 4676 77598
rect 4620 76468 4676 77532
rect 4732 77364 4788 77374
rect 4732 76690 4788 77308
rect 4732 76638 4734 76690
rect 4786 76638 4788 76690
rect 4732 76626 4788 76638
rect 4732 76468 4788 76478
rect 4620 76466 4788 76468
rect 4620 76414 4734 76466
rect 4786 76414 4788 76466
rect 4620 76412 4788 76414
rect 4732 76402 4788 76412
rect 4508 76290 4564 76300
rect 4620 76244 4676 76282
rect 4620 76178 4676 76188
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4284 75684 4340 75694
rect 4508 75684 4564 75722
rect 4284 75682 4452 75684
rect 4284 75630 4286 75682
rect 4338 75630 4452 75682
rect 4284 75628 4452 75630
rect 4284 75618 4340 75628
rect 3948 75506 4004 75516
rect 4060 75516 4228 75572
rect 4396 75572 4452 75628
rect 4508 75618 4564 75628
rect 3836 75394 3892 75404
rect 4060 75236 4116 75516
rect 4396 75506 4452 75516
rect 4732 75572 4788 75582
rect 4732 75478 4788 75516
rect 3612 75180 3780 75236
rect 3836 75180 4116 75236
rect 4508 75458 4564 75470
rect 4508 75406 4510 75458
rect 4562 75406 4564 75458
rect 3500 74004 3556 74042
rect 3500 73938 3556 73948
rect 3388 73490 3444 73500
rect 3276 73218 3332 73230
rect 3276 73166 3278 73218
rect 3330 73166 3332 73218
rect 3276 72436 3332 73166
rect 3388 72770 3444 72782
rect 3388 72718 3390 72770
rect 3442 72718 3444 72770
rect 3388 72658 3444 72718
rect 3388 72606 3390 72658
rect 3442 72606 3444 72658
rect 3388 72594 3444 72606
rect 3276 72370 3332 72380
rect 3612 72212 3668 75180
rect 3836 75124 3892 75180
rect 3724 75068 3892 75124
rect 3724 73444 3780 75068
rect 4060 75012 4116 75022
rect 3836 74786 3892 74798
rect 3836 74734 3838 74786
rect 3890 74734 3892 74786
rect 3836 73892 3892 74734
rect 3948 74004 4004 74042
rect 3948 73938 4004 73948
rect 3836 73826 3892 73836
rect 3724 73388 3892 73444
rect 3724 73220 3780 73230
rect 3724 73126 3780 73164
rect 3836 72770 3892 73388
rect 4060 73220 4116 74956
rect 4172 74788 4228 74798
rect 4172 73442 4228 74732
rect 4508 74788 4564 75406
rect 4508 74722 4564 74732
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4844 74226 4900 78428
rect 4956 77364 5012 79436
rect 7168 79200 7280 80000
rect 10892 79604 10948 79614
rect 8316 79380 8372 79390
rect 7196 79044 7252 79200
rect 7196 78988 7476 79044
rect 4956 77298 5012 77308
rect 5852 78932 5908 78942
rect 5852 76690 5908 78876
rect 7084 77700 7140 77710
rect 7084 77606 7140 77644
rect 5852 76638 5854 76690
rect 5906 76638 5908 76690
rect 5852 76626 5908 76638
rect 6636 76804 6692 76814
rect 6300 76468 6356 76478
rect 6300 76374 6356 76412
rect 6636 76466 6692 76748
rect 7420 76580 7476 78988
rect 7644 78260 7700 78270
rect 7532 76580 7588 76590
rect 7420 76578 7588 76580
rect 7420 76526 7534 76578
rect 7586 76526 7588 76578
rect 7420 76524 7588 76526
rect 6636 76414 6638 76466
rect 6690 76414 6692 76466
rect 6636 76356 6692 76414
rect 6860 76466 6916 76478
rect 6860 76414 6862 76466
rect 6914 76414 6916 76466
rect 6636 76290 6692 76300
rect 6748 76354 6804 76366
rect 6748 76302 6750 76354
rect 6802 76302 6804 76354
rect 5628 76244 5684 76254
rect 5404 75908 5460 75918
rect 4956 75570 5012 75582
rect 4956 75518 4958 75570
rect 5010 75518 5012 75570
rect 4956 74900 5012 75518
rect 4956 74834 5012 74844
rect 5180 75012 5236 75022
rect 4844 74174 4846 74226
rect 4898 74174 4900 74226
rect 4844 74162 4900 74174
rect 4956 74340 5012 74350
rect 4396 74116 4452 74126
rect 4396 74022 4452 74060
rect 4732 74116 4788 74154
rect 4732 74050 4788 74060
rect 4956 74114 5012 74284
rect 4956 74062 4958 74114
rect 5010 74062 5012 74114
rect 4956 74050 5012 74062
rect 4172 73390 4174 73442
rect 4226 73390 4228 73442
rect 4172 73378 4228 73390
rect 4844 73780 4900 73790
rect 4508 73330 4564 73342
rect 4508 73278 4510 73330
rect 4562 73278 4564 73330
rect 4284 73220 4340 73230
rect 4060 73218 4340 73220
rect 4060 73166 4286 73218
rect 4338 73166 4340 73218
rect 4060 73164 4340 73166
rect 4284 73154 4340 73164
rect 4508 73108 4564 73278
rect 4508 73042 4564 73052
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 3836 72718 3838 72770
rect 3890 72718 3892 72770
rect 3836 72706 3892 72718
rect 4284 72772 4340 72782
rect 3500 72156 3668 72212
rect 3724 72660 3780 72670
rect 3388 71764 3444 71802
rect 3388 71698 3444 71708
rect 3388 71540 3444 71550
rect 3388 70084 3444 71484
rect 3500 71090 3556 72156
rect 3724 72100 3780 72604
rect 4284 72658 4340 72716
rect 4284 72606 4286 72658
rect 4338 72606 4340 72658
rect 4284 72594 4340 72606
rect 4508 72770 4564 72782
rect 4844 72772 4900 73724
rect 5180 73332 5236 74956
rect 5292 74900 5348 74910
rect 5292 74116 5348 74844
rect 5292 74050 5348 74060
rect 5180 73238 5236 73276
rect 5404 73330 5460 75852
rect 5404 73278 5406 73330
rect 5458 73278 5460 73330
rect 5404 73266 5460 73278
rect 4508 72718 4510 72770
rect 4562 72718 4564 72770
rect 3836 72548 3892 72558
rect 3836 72454 3892 72492
rect 3500 71038 3502 71090
rect 3554 71038 3556 71090
rect 3500 71026 3556 71038
rect 3612 72044 3780 72100
rect 3388 70082 3556 70084
rect 3388 70030 3390 70082
rect 3442 70030 3556 70082
rect 3388 70028 3556 70030
rect 3388 70018 3444 70028
rect 3164 69804 3332 69860
rect 3164 69524 3220 69534
rect 3164 69430 3220 69468
rect 3276 69300 3332 69804
rect 2940 68674 2996 68684
rect 3052 69244 3332 69300
rect 2940 68514 2996 68526
rect 2940 68462 2942 68514
rect 2994 68462 2996 68514
rect 2828 67844 2884 67854
rect 2828 67750 2884 67788
rect 2716 67116 2884 67172
rect 2604 67106 2660 67116
rect 2380 66948 2436 66958
rect 2380 66946 2548 66948
rect 2380 66894 2382 66946
rect 2434 66894 2548 66946
rect 2380 66892 2548 66894
rect 2380 66882 2436 66892
rect 2156 66334 2158 66386
rect 2210 66334 2212 66386
rect 2156 64148 2212 66334
rect 2268 65492 2324 65502
rect 2268 65398 2324 65436
rect 2380 64820 2436 64830
rect 1932 64082 1988 64092
rect 2156 64082 2212 64092
rect 2268 64708 2324 64718
rect 1820 63970 1876 63980
rect 1708 63646 1710 63698
rect 1762 63646 1764 63698
rect 1708 63634 1764 63646
rect 1932 63812 1988 63822
rect 1932 63250 1988 63756
rect 1932 63198 1934 63250
rect 1986 63198 1988 63250
rect 1932 63186 1988 63198
rect 1932 62580 1988 62590
rect 2268 62580 2324 64652
rect 2380 64260 2436 64764
rect 2380 64194 2436 64204
rect 2380 63924 2436 63934
rect 2380 63830 2436 63868
rect 2492 63588 2548 66892
rect 2716 66946 2772 66958
rect 2716 66894 2718 66946
rect 2770 66894 2772 66946
rect 2716 66500 2772 66894
rect 2716 66434 2772 66444
rect 2604 66388 2660 66398
rect 2604 66294 2660 66332
rect 2716 65378 2772 65390
rect 2716 65326 2718 65378
rect 2770 65326 2772 65378
rect 2716 65156 2772 65326
rect 2716 65090 2772 65100
rect 2492 63522 2548 63532
rect 2604 64930 2660 64942
rect 2604 64878 2606 64930
rect 2658 64878 2660 64930
rect 2604 64148 2660 64878
rect 2828 64820 2884 67116
rect 2940 66948 2996 68462
rect 2940 66882 2996 66892
rect 2828 64754 2884 64764
rect 2940 66500 2996 66510
rect 2828 64596 2884 64606
rect 2828 64502 2884 64540
rect 2716 64148 2772 64158
rect 2604 64146 2772 64148
rect 2604 64094 2718 64146
rect 2770 64094 2772 64146
rect 2604 64092 2772 64094
rect 2492 63362 2548 63374
rect 2492 63310 2494 63362
rect 2546 63310 2548 63362
rect 2380 63140 2436 63150
rect 2380 63046 2436 63084
rect 1932 62578 2324 62580
rect 1932 62526 1934 62578
rect 1986 62526 2324 62578
rect 1932 62524 2324 62526
rect 2380 62580 2436 62590
rect 2492 62580 2548 63310
rect 2604 62692 2660 64092
rect 2716 64082 2772 64092
rect 2940 63812 2996 66444
rect 3052 65716 3108 69244
rect 3388 68740 3444 68750
rect 3388 68514 3444 68684
rect 3388 68462 3390 68514
rect 3442 68462 3444 68514
rect 3164 68068 3220 68078
rect 3164 67396 3220 68012
rect 3388 67956 3444 68462
rect 3388 67890 3444 67900
rect 3276 67732 3332 67742
rect 3276 67638 3332 67676
rect 3164 67330 3220 67340
rect 3164 67172 3220 67182
rect 3164 66500 3220 67116
rect 3500 67060 3556 70028
rect 3612 68740 3668 72044
rect 3724 71876 3780 71886
rect 3724 69860 3780 71820
rect 3836 71764 3892 71774
rect 3836 71670 3892 71708
rect 4284 71650 4340 71662
rect 4284 71598 4286 71650
rect 4338 71598 4340 71650
rect 4284 71540 4340 71598
rect 4060 71484 4340 71540
rect 4508 71540 4564 72718
rect 4732 72716 4900 72772
rect 4956 73220 5012 73230
rect 4732 72434 4788 72716
rect 4732 72382 4734 72434
rect 4786 72382 4788 72434
rect 4732 71652 4788 72382
rect 4844 72322 4900 72334
rect 4844 72270 4846 72322
rect 4898 72270 4900 72322
rect 4844 72212 4900 72270
rect 4844 72146 4900 72156
rect 4732 71586 4788 71596
rect 4844 71650 4900 71662
rect 4844 71598 4846 71650
rect 4898 71598 4900 71650
rect 3948 71092 4004 71102
rect 3948 70998 4004 71036
rect 3836 70196 3892 70206
rect 3836 70102 3892 70140
rect 3724 69804 3892 69860
rect 3724 69412 3780 69422
rect 3724 69318 3780 69356
rect 3612 68674 3668 68684
rect 3724 68852 3780 68862
rect 3724 68404 3780 68796
rect 3836 68740 3892 69804
rect 3836 68674 3892 68684
rect 3612 68348 3780 68404
rect 3836 68514 3892 68526
rect 3836 68462 3838 68514
rect 3890 68462 3892 68514
rect 3612 67282 3668 68348
rect 3612 67230 3614 67282
rect 3666 67230 3668 67282
rect 3612 67218 3668 67230
rect 3724 68180 3780 68190
rect 3724 67954 3780 68124
rect 3724 67902 3726 67954
rect 3778 67902 3780 67954
rect 3724 67172 3780 67902
rect 3836 67284 3892 68462
rect 3836 67218 3892 67228
rect 3724 67106 3780 67116
rect 3164 66434 3220 66444
rect 3276 67004 3556 67060
rect 3052 65650 3108 65660
rect 3164 66274 3220 66286
rect 3164 66222 3166 66274
rect 3218 66222 3220 66274
rect 3052 65378 3108 65390
rect 3052 65326 3054 65378
rect 3106 65326 3108 65378
rect 3052 65156 3108 65326
rect 3052 65090 3108 65100
rect 3164 64932 3220 66222
rect 3276 65940 3332 67004
rect 3724 66948 3780 66958
rect 3388 66834 3444 66846
rect 3388 66782 3390 66834
rect 3442 66782 3444 66834
rect 3388 66162 3444 66782
rect 3388 66110 3390 66162
rect 3442 66110 3444 66162
rect 3388 66098 3444 66110
rect 3276 65884 3444 65940
rect 3164 64866 3220 64876
rect 3164 64708 3220 64718
rect 3388 64708 3444 65884
rect 3612 65378 3668 65390
rect 3612 65326 3614 65378
rect 3666 65326 3668 65378
rect 3612 64932 3668 65326
rect 3164 64614 3220 64652
rect 3276 64652 3444 64708
rect 3500 64930 3668 64932
rect 3500 64878 3614 64930
rect 3666 64878 3668 64930
rect 3500 64876 3668 64878
rect 3164 63812 3220 63850
rect 2940 63756 3164 63812
rect 3164 63746 3220 63756
rect 2828 63698 2884 63710
rect 2828 63646 2830 63698
rect 2882 63646 2884 63698
rect 2716 63476 2772 63486
rect 2716 63250 2772 63420
rect 2716 63198 2718 63250
rect 2770 63198 2772 63250
rect 2716 62804 2772 63198
rect 2716 62738 2772 62748
rect 2604 62626 2660 62636
rect 2380 62578 2548 62580
rect 2380 62526 2382 62578
rect 2434 62526 2548 62578
rect 2380 62524 2548 62526
rect 2716 62580 2772 62590
rect 2828 62580 2884 63646
rect 3164 63588 3220 63598
rect 3164 63250 3220 63532
rect 3276 63362 3332 64652
rect 3276 63310 3278 63362
rect 3330 63310 3332 63362
rect 3276 63298 3332 63310
rect 3388 64484 3444 64494
rect 3164 63198 3166 63250
rect 3218 63198 3220 63250
rect 3164 62804 3220 63198
rect 3164 62738 3220 62748
rect 2716 62578 2884 62580
rect 2716 62526 2718 62578
rect 2770 62526 2884 62578
rect 2716 62524 2884 62526
rect 3276 62692 3332 62702
rect 3276 62578 3332 62636
rect 3276 62526 3278 62578
rect 3330 62526 3332 62578
rect 1932 62514 1988 62524
rect 1932 61348 1988 61358
rect 1932 61254 1988 61292
rect 1932 61012 1988 61022
rect 1932 60918 1988 60956
rect 2044 60116 2100 62524
rect 2380 62188 2436 62524
rect 2716 62468 2772 62524
rect 3276 62514 3332 62526
rect 2268 62132 2436 62188
rect 2492 62412 2772 62468
rect 2268 61012 2324 62132
rect 2492 61796 2548 62412
rect 2828 62356 2884 62366
rect 2716 62300 2828 62356
rect 2492 61730 2548 61740
rect 2604 62244 2660 62254
rect 2380 61684 2436 61694
rect 2380 61590 2436 61628
rect 2604 61572 2660 62188
rect 2492 61516 2660 61572
rect 2716 61682 2772 62300
rect 2828 62290 2884 62300
rect 3052 62356 3108 62366
rect 2716 61630 2718 61682
rect 2770 61630 2772 61682
rect 2716 61572 2772 61630
rect 2380 61012 2436 61022
rect 2268 61010 2436 61012
rect 2268 60958 2382 61010
rect 2434 60958 2436 61010
rect 2268 60956 2436 60958
rect 2380 60946 2436 60956
rect 2156 60116 2212 60126
rect 2044 60114 2212 60116
rect 2044 60062 2158 60114
rect 2210 60062 2212 60114
rect 2044 60060 2212 60062
rect 1596 60050 1652 60060
rect 2156 60050 2212 60060
rect 2492 59892 2548 61516
rect 2604 60228 2660 60238
rect 2604 60114 2660 60172
rect 2604 60062 2606 60114
rect 2658 60062 2660 60114
rect 2604 60050 2660 60062
rect 2492 59826 2548 59836
rect 2716 50036 2772 61516
rect 2828 62188 2884 62198
rect 3052 62188 3108 62300
rect 2828 61010 2884 62132
rect 2828 60958 2830 61010
rect 2882 60958 2884 61010
rect 2828 54516 2884 60958
rect 2940 62132 3108 62188
rect 3388 62132 3444 64428
rect 3500 63812 3556 64876
rect 3612 64866 3668 64876
rect 3612 64708 3668 64718
rect 3612 64036 3668 64652
rect 3724 64260 3780 66892
rect 4060 66612 4116 71484
rect 4508 71474 4564 71484
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4172 71204 4228 71214
rect 4172 69522 4228 71148
rect 4844 71204 4900 71598
rect 4844 71138 4900 71148
rect 4620 71092 4676 71102
rect 4508 71036 4620 71092
rect 4396 70980 4452 70990
rect 4396 70886 4452 70924
rect 4508 70756 4564 71036
rect 4620 70998 4676 71036
rect 4956 71092 5012 73164
rect 5068 73106 5124 73118
rect 5068 73054 5070 73106
rect 5122 73054 5124 73106
rect 5068 72548 5124 73054
rect 5516 73108 5572 73118
rect 5516 73014 5572 73052
rect 5292 72548 5348 72558
rect 5068 72492 5236 72548
rect 5068 72322 5124 72334
rect 5068 72270 5070 72322
rect 5122 72270 5124 72322
rect 5068 71876 5124 72270
rect 5068 71810 5124 71820
rect 4956 71026 5012 71036
rect 4172 69470 4174 69522
rect 4226 69470 4228 69522
rect 4172 69458 4228 69470
rect 4284 70700 4564 70756
rect 4844 70980 4900 70990
rect 4284 69300 4340 70700
rect 4396 70532 4452 70542
rect 4396 70418 4452 70476
rect 4396 70366 4398 70418
rect 4450 70366 4452 70418
rect 4396 70354 4452 70366
rect 4844 70196 4900 70924
rect 4956 70756 5012 70766
rect 4956 70662 5012 70700
rect 5180 70420 5236 72492
rect 5068 70364 5236 70420
rect 4844 70140 5012 70196
rect 4732 70084 4788 70094
rect 4732 70082 4900 70084
rect 4732 70030 4734 70082
rect 4786 70030 4900 70082
rect 4732 70028 4900 70030
rect 4732 70018 4788 70028
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 4508 69524 4564 69534
rect 4508 69430 4564 69468
rect 4284 69234 4340 69244
rect 4844 69188 4900 70028
rect 4396 68740 4452 68750
rect 4396 68646 4452 68684
rect 4844 68628 4900 69132
rect 4844 68562 4900 68572
rect 4956 69522 5012 70140
rect 5068 69748 5124 70364
rect 5180 70194 5236 70206
rect 5180 70142 5182 70194
rect 5234 70142 5236 70194
rect 5180 70084 5236 70142
rect 5180 70018 5236 70028
rect 5068 69682 5124 69692
rect 4956 69470 4958 69522
rect 5010 69470 5012 69522
rect 4284 68402 4340 68414
rect 4284 68350 4286 68402
rect 4338 68350 4340 68402
rect 4284 68292 4340 68350
rect 4284 68226 4340 68236
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4844 68180 4900 68190
rect 4844 68068 4900 68124
rect 4508 68012 4900 68068
rect 4172 67844 4228 67854
rect 4508 67844 4564 68012
rect 4172 67842 4564 67844
rect 4172 67790 4174 67842
rect 4226 67790 4564 67842
rect 4172 67788 4564 67790
rect 4620 67844 4676 67854
rect 4956 67844 5012 69470
rect 5068 69188 5124 69198
rect 5068 68850 5124 69132
rect 5068 68798 5070 68850
rect 5122 68798 5124 68850
rect 5068 68786 5124 68798
rect 4172 67778 4228 67788
rect 4620 67750 4676 67788
rect 4844 67788 5012 67844
rect 5068 68628 5124 68638
rect 5292 68628 5348 72492
rect 5404 72100 5460 72110
rect 5404 71874 5460 72044
rect 5628 71986 5684 76188
rect 6300 76244 6356 76254
rect 5964 75908 6020 75918
rect 5740 74228 5796 74238
rect 5740 72100 5796 74172
rect 5964 74226 6020 75852
rect 6076 75794 6132 75806
rect 6076 75742 6078 75794
rect 6130 75742 6132 75794
rect 6076 75012 6132 75742
rect 6076 74956 6244 75012
rect 6076 74786 6132 74798
rect 6076 74734 6078 74786
rect 6130 74734 6132 74786
rect 6076 74676 6132 74734
rect 6076 74610 6132 74620
rect 5964 74174 5966 74226
rect 6018 74174 6020 74226
rect 5964 74162 6020 74174
rect 6188 73556 6244 74956
rect 6188 73490 6244 73500
rect 6188 73332 6244 73342
rect 6300 73332 6356 76188
rect 6748 76132 6804 76302
rect 6748 76066 6804 76076
rect 6860 75908 6916 76414
rect 6524 75852 6916 75908
rect 7308 76468 7364 76478
rect 6412 73892 6468 73902
rect 6412 73798 6468 73836
rect 6244 73276 6356 73332
rect 6412 73332 6468 73342
rect 6188 73238 6244 73276
rect 6412 73238 6468 73276
rect 5740 72034 5796 72044
rect 5852 73108 5908 73118
rect 5852 72436 5908 73052
rect 6300 72772 6356 72782
rect 6300 72678 6356 72716
rect 6188 72548 6244 72558
rect 5964 72436 6020 72446
rect 5852 72434 6020 72436
rect 5852 72382 5966 72434
rect 6018 72382 6020 72434
rect 5852 72380 6020 72382
rect 5628 71934 5630 71986
rect 5682 71934 5684 71986
rect 5628 71922 5684 71934
rect 5404 71822 5406 71874
rect 5458 71822 5460 71874
rect 5404 70756 5460 71822
rect 5740 71876 5796 71886
rect 5740 71782 5796 71820
rect 5404 70690 5460 70700
rect 5516 71540 5572 71550
rect 4284 67172 4340 67182
rect 4172 66948 4228 66958
rect 4172 66854 4228 66892
rect 4060 66556 4228 66612
rect 4060 66388 4116 66398
rect 3836 66332 4060 66388
rect 3836 65492 3892 66332
rect 4060 66294 4116 66332
rect 3836 65426 3892 65436
rect 4060 65492 4116 65502
rect 4060 65398 4116 65436
rect 4060 64484 4116 64494
rect 4060 64390 4116 64428
rect 3724 64204 4116 64260
rect 3612 63970 3668 63980
rect 3948 64036 4004 64046
rect 3724 63924 3780 63934
rect 3724 63830 3780 63868
rect 3500 63756 3668 63812
rect 3612 63588 3668 63756
rect 3612 63532 3780 63588
rect 2940 57764 2996 62132
rect 3276 62076 3444 62132
rect 3500 63476 3556 63486
rect 3164 61796 3220 61806
rect 3164 61682 3220 61740
rect 3164 61630 3166 61682
rect 3218 61630 3220 61682
rect 3164 61618 3220 61630
rect 3164 61236 3220 61246
rect 3164 61010 3220 61180
rect 3164 60958 3166 61010
rect 3218 60958 3220 61010
rect 3164 60946 3220 60958
rect 3276 61012 3332 62076
rect 3276 60946 3332 60956
rect 3388 61794 3444 61806
rect 3388 61742 3390 61794
rect 3442 61742 3444 61794
rect 3052 60116 3108 60126
rect 3052 59332 3108 60060
rect 3388 60114 3444 61742
rect 3500 60226 3556 63420
rect 3612 63364 3668 63374
rect 3612 63250 3668 63308
rect 3612 63198 3614 63250
rect 3666 63198 3668 63250
rect 3612 63186 3668 63198
rect 3612 62580 3668 62590
rect 3724 62580 3780 63532
rect 3612 62578 3780 62580
rect 3612 62526 3614 62578
rect 3666 62526 3780 62578
rect 3612 62524 3780 62526
rect 3612 62514 3668 62524
rect 3724 61796 3780 62524
rect 3724 61730 3780 61740
rect 3612 61348 3668 61358
rect 3612 61254 3668 61292
rect 3500 60174 3502 60226
rect 3554 60174 3556 60226
rect 3500 60162 3556 60174
rect 3724 60788 3780 60798
rect 3724 60674 3780 60732
rect 3724 60622 3726 60674
rect 3778 60622 3780 60674
rect 3388 60062 3390 60114
rect 3442 60062 3444 60114
rect 3388 60050 3444 60062
rect 3052 59266 3108 59276
rect 3388 59444 3444 59454
rect 3388 59106 3444 59388
rect 3388 59054 3390 59106
rect 3442 59054 3444 59106
rect 3388 57876 3444 59054
rect 3724 58660 3780 60622
rect 3948 60114 4004 63980
rect 4060 63810 4116 64204
rect 4060 63758 4062 63810
rect 4114 63758 4116 63810
rect 4060 63698 4116 63758
rect 4060 63646 4062 63698
rect 4114 63646 4116 63698
rect 4060 61794 4116 63646
rect 4172 63700 4228 66556
rect 4284 66388 4340 67116
rect 4508 67172 4564 67182
rect 4508 66836 4564 67116
rect 4844 67170 4900 67788
rect 4844 67118 4846 67170
rect 4898 67118 4900 67170
rect 4844 67106 4900 67118
rect 4956 67618 5012 67630
rect 4956 67566 4958 67618
rect 5010 67566 5012 67618
rect 4956 67172 5012 67566
rect 4956 67106 5012 67116
rect 4620 67060 4676 67070
rect 4620 66966 4676 67004
rect 4956 66946 5012 66958
rect 4956 66894 4958 66946
rect 5010 66894 5012 66946
rect 4508 66780 4900 66836
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4508 66500 4564 66510
rect 4844 66500 4900 66780
rect 4956 66612 5012 66894
rect 5068 66948 5124 68572
rect 5180 68572 5348 68628
rect 5404 69524 5460 69534
rect 5404 68964 5460 69468
rect 5180 68514 5236 68572
rect 5180 68462 5182 68514
rect 5234 68462 5236 68514
rect 5180 68450 5236 68462
rect 5292 68404 5348 68414
rect 5292 68310 5348 68348
rect 5404 67170 5460 68908
rect 5516 68066 5572 71484
rect 5852 71316 5908 72380
rect 5964 72370 6020 72380
rect 6188 72324 6244 72492
rect 6188 72230 6244 72268
rect 6300 72212 6356 72222
rect 6188 72100 6244 72110
rect 5964 71764 6020 71774
rect 5964 71670 6020 71708
rect 5628 71260 5908 71316
rect 5964 71428 6020 71438
rect 5628 71202 5684 71260
rect 5628 71150 5630 71202
rect 5682 71150 5684 71202
rect 5628 71138 5684 71150
rect 5964 70978 6020 71372
rect 5964 70926 5966 70978
rect 6018 70926 6020 70978
rect 5964 70914 6020 70926
rect 5852 70756 5908 70766
rect 6188 70756 6244 72044
rect 6300 71316 6356 72156
rect 6524 71874 6580 75852
rect 6860 75684 6916 75694
rect 6860 74898 6916 75628
rect 6860 74846 6862 74898
rect 6914 74846 6916 74898
rect 6860 74834 6916 74846
rect 7196 75572 7252 75582
rect 7084 74452 7140 74462
rect 7084 74338 7140 74396
rect 7084 74286 7086 74338
rect 7138 74286 7140 74338
rect 7084 74274 7140 74286
rect 6972 74114 7028 74126
rect 6972 74062 6974 74114
rect 7026 74062 7028 74114
rect 6972 74004 7028 74062
rect 6972 73938 7028 73948
rect 7196 74004 7252 75516
rect 6748 73892 6804 73902
rect 6748 73442 6804 73836
rect 6748 73390 6750 73442
rect 6802 73390 6804 73442
rect 6748 73378 6804 73390
rect 6972 73556 7028 73566
rect 6636 73218 6692 73230
rect 6636 73166 6638 73218
rect 6690 73166 6692 73218
rect 6636 72660 6692 73166
rect 6636 72594 6692 72604
rect 6860 72548 6916 72558
rect 6860 72454 6916 72492
rect 6524 71822 6526 71874
rect 6578 71822 6580 71874
rect 6524 71810 6580 71822
rect 6300 70978 6356 71260
rect 6300 70926 6302 70978
rect 6354 70926 6356 70978
rect 6300 70914 6356 70926
rect 6412 71092 6468 71102
rect 6412 70978 6468 71036
rect 6412 70926 6414 70978
rect 6466 70926 6468 70978
rect 6412 70914 6468 70926
rect 6524 70980 6580 70990
rect 6524 70886 6580 70924
rect 6412 70756 6468 70766
rect 6188 70700 6356 70756
rect 5628 70420 5684 70430
rect 5628 70326 5684 70364
rect 5852 70418 5908 70700
rect 6076 70644 6132 70654
rect 5852 70366 5854 70418
rect 5906 70366 5908 70418
rect 5852 70354 5908 70366
rect 5964 70532 6132 70588
rect 5740 70082 5796 70094
rect 5740 70030 5742 70082
rect 5794 70030 5796 70082
rect 5516 68014 5518 68066
rect 5570 68014 5572 68066
rect 5516 68002 5572 68014
rect 5628 69748 5684 69758
rect 5628 67844 5684 69692
rect 5740 69300 5796 70030
rect 5852 69636 5908 69646
rect 5852 69542 5908 69580
rect 5740 69234 5796 69244
rect 5964 69410 6020 70532
rect 6300 70420 6356 70700
rect 6300 70354 6356 70364
rect 6188 70308 6244 70318
rect 6188 69634 6244 70252
rect 6188 69582 6190 69634
rect 6242 69582 6244 69634
rect 6188 69570 6244 69582
rect 6300 69636 6356 69646
rect 6300 69542 6356 69580
rect 5964 69358 5966 69410
rect 6018 69358 6020 69410
rect 5964 68740 6020 69358
rect 5964 68674 6020 68684
rect 6076 69300 6132 69310
rect 6076 68514 6132 69244
rect 6076 68462 6078 68514
rect 6130 68462 6132 68514
rect 6076 68450 6132 68462
rect 5740 68068 5796 68078
rect 5740 68066 6020 68068
rect 5740 68014 5742 68066
rect 5794 68014 6020 68066
rect 5740 68012 6020 68014
rect 5740 68002 5796 68012
rect 5404 67118 5406 67170
rect 5458 67118 5460 67170
rect 5404 67106 5460 67118
rect 5516 67788 5684 67844
rect 5964 67842 6020 68012
rect 5964 67790 5966 67842
rect 6018 67790 6020 67842
rect 5180 66948 5236 66958
rect 5068 66892 5180 66948
rect 4956 66546 5012 66556
rect 4284 66332 4452 66388
rect 4284 66164 4340 66174
rect 4284 64820 4340 66108
rect 4396 66052 4452 66332
rect 4396 65986 4452 65996
rect 4508 65828 4564 66444
rect 4620 66444 4900 66500
rect 4620 66386 4676 66444
rect 4620 66334 4622 66386
rect 4674 66334 4676 66386
rect 4620 66322 4676 66334
rect 5068 66050 5124 66062
rect 5068 65998 5070 66050
rect 5122 65998 5124 66050
rect 4508 65762 4564 65772
rect 4620 65940 4676 65950
rect 4508 65378 4564 65390
rect 4508 65326 4510 65378
rect 4562 65326 4564 65378
rect 4508 65266 4564 65326
rect 4620 65380 4676 65884
rect 5068 65828 5124 65998
rect 5068 65762 5124 65772
rect 4844 65604 4900 65614
rect 5180 65604 5236 66892
rect 5516 65828 5572 67788
rect 5852 66948 5908 66958
rect 5852 66854 5908 66892
rect 5964 66498 6020 67790
rect 5964 66446 5966 66498
rect 6018 66446 6020 66498
rect 5516 65762 5572 65772
rect 5740 66050 5796 66062
rect 5740 65998 5742 66050
rect 5794 65998 5796 66050
rect 5628 65716 5684 65726
rect 4900 65548 5236 65604
rect 5404 65604 5460 65614
rect 4844 65472 4900 65548
rect 5404 65490 5460 65548
rect 5404 65438 5406 65490
rect 5458 65438 5460 65490
rect 5404 65426 5460 65438
rect 4620 65324 5012 65380
rect 4508 65214 4510 65266
rect 4562 65214 4564 65266
rect 4508 65202 4564 65214
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4956 65044 5012 65324
rect 4956 64978 5012 64988
rect 5180 65266 5236 65278
rect 5180 65214 5182 65266
rect 5234 65214 5236 65266
rect 4956 64820 5012 64830
rect 4284 64764 4676 64820
rect 4508 64596 4564 64606
rect 4508 64502 4564 64540
rect 4620 64146 4676 64764
rect 4956 64726 5012 64764
rect 4844 64706 4900 64718
rect 4844 64654 4846 64706
rect 4898 64654 4900 64706
rect 4844 64484 4900 64654
rect 5180 64596 5236 65214
rect 5516 65268 5572 65278
rect 5516 65174 5572 65212
rect 5180 64530 5236 64540
rect 4844 64418 4900 64428
rect 4620 64094 4622 64146
rect 4674 64094 4676 64146
rect 4620 64082 4676 64094
rect 5516 64148 5572 64158
rect 5628 64148 5684 65660
rect 5740 65380 5796 65998
rect 5740 65314 5796 65324
rect 5852 65716 5908 65726
rect 5572 64092 5684 64148
rect 5852 64146 5908 65660
rect 5852 64094 5854 64146
rect 5906 64094 5908 64146
rect 5516 64054 5572 64092
rect 4172 63634 4228 63644
rect 4844 63812 4900 63822
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4172 63364 4228 63374
rect 4172 63250 4228 63308
rect 4172 63198 4174 63250
rect 4226 63198 4228 63250
rect 4172 63186 4228 63198
rect 4508 63362 4564 63374
rect 4508 63310 4510 63362
rect 4562 63310 4564 63362
rect 4508 62804 4564 63310
rect 4620 63252 4676 63262
rect 4620 63158 4676 63196
rect 4508 62578 4564 62748
rect 4508 62526 4510 62578
rect 4562 62526 4564 62578
rect 4508 62514 4564 62526
rect 4844 62916 4900 63756
rect 4956 63812 5012 63822
rect 4956 63810 5124 63812
rect 4956 63758 4958 63810
rect 5010 63758 5124 63810
rect 4956 63756 5124 63758
rect 4956 63746 5012 63756
rect 4956 62916 5012 62926
rect 4844 62914 5012 62916
rect 4844 62862 4958 62914
rect 5010 62862 5012 62914
rect 4844 62860 5012 62862
rect 4844 62354 4900 62860
rect 4956 62850 5012 62860
rect 4844 62302 4846 62354
rect 4898 62302 4900 62354
rect 4844 62290 4900 62302
rect 4956 62356 5012 62366
rect 4172 62244 4228 62282
rect 4956 62262 5012 62300
rect 4172 62178 4228 62188
rect 4844 62132 4900 62142
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 4060 61742 4062 61794
rect 4114 61742 4116 61794
rect 4060 61730 4116 61742
rect 4172 61684 4228 61694
rect 4060 61572 4116 61582
rect 4060 61478 4116 61516
rect 4172 61010 4228 61628
rect 4508 61684 4564 61694
rect 4508 61590 4564 61628
rect 4172 60958 4174 61010
rect 4226 60958 4228 61010
rect 4172 60946 4228 60958
rect 4396 61236 4452 61246
rect 4396 60788 4452 61180
rect 4172 60732 4452 60788
rect 3948 60062 3950 60114
rect 4002 60062 4004 60114
rect 3948 60050 4004 60062
rect 4060 60676 4116 60686
rect 3948 59444 4004 59454
rect 4060 59444 4116 60620
rect 3948 59442 4116 59444
rect 3948 59390 3950 59442
rect 4002 59390 4116 59442
rect 3948 59388 4116 59390
rect 3948 59378 4004 59388
rect 3724 58594 3780 58604
rect 4172 58996 4228 60732
rect 4508 60676 4564 60686
rect 4844 60676 4900 62076
rect 4956 61684 5012 61694
rect 5068 61684 5124 63756
rect 5852 63252 5908 64094
rect 5852 63186 5908 63196
rect 5964 64820 6020 66446
rect 6076 67618 6132 67630
rect 6076 67566 6078 67618
rect 6130 67566 6132 67618
rect 6076 67172 6132 67566
rect 6300 67618 6356 67630
rect 6300 67566 6302 67618
rect 6354 67566 6356 67618
rect 6300 67508 6356 67566
rect 6300 67442 6356 67452
rect 6076 65716 6132 67116
rect 6076 65650 6132 65660
rect 6188 67284 6244 67294
rect 6412 67284 6468 70700
rect 6748 70644 6804 70654
rect 6636 70532 6804 70588
rect 6636 69748 6692 70532
rect 6748 70420 6804 70430
rect 6748 70326 6804 70364
rect 6860 70306 6916 70318
rect 6860 70254 6862 70306
rect 6914 70254 6916 70306
rect 6860 70196 6916 70254
rect 6524 69692 6636 69748
rect 6524 69188 6580 69692
rect 6636 69682 6692 69692
rect 6748 70140 6916 70196
rect 6524 69122 6580 69132
rect 6636 69300 6692 69310
rect 6076 64820 6132 64830
rect 6020 64818 6132 64820
rect 6020 64766 6078 64818
rect 6130 64766 6132 64818
rect 6020 64764 6132 64766
rect 5516 62580 5572 62590
rect 5964 62580 6020 64764
rect 6076 64754 6132 64764
rect 5516 62578 6020 62580
rect 5516 62526 5518 62578
rect 5570 62526 5966 62578
rect 6018 62526 6020 62578
rect 5516 62524 6020 62526
rect 5516 62514 5572 62524
rect 5964 62514 6020 62524
rect 6076 62914 6132 62926
rect 6076 62862 6078 62914
rect 6130 62862 6132 62914
rect 6076 62132 6132 62862
rect 6188 62188 6244 67228
rect 6300 67228 6468 67284
rect 6524 67620 6580 67630
rect 6300 66386 6356 67228
rect 6524 66948 6580 67564
rect 6636 67282 6692 69244
rect 6636 67230 6638 67282
rect 6690 67230 6692 67282
rect 6636 67172 6692 67230
rect 6636 67106 6692 67116
rect 6636 66948 6692 66958
rect 6524 66946 6692 66948
rect 6524 66894 6638 66946
rect 6690 66894 6692 66946
rect 6524 66892 6692 66894
rect 6412 66834 6468 66846
rect 6412 66782 6414 66834
rect 6466 66782 6468 66834
rect 6412 66498 6468 66782
rect 6412 66446 6414 66498
rect 6466 66446 6468 66498
rect 6412 66434 6468 66446
rect 6300 66334 6302 66386
rect 6354 66334 6356 66386
rect 6300 66322 6356 66334
rect 6524 65716 6580 65726
rect 6300 65378 6356 65390
rect 6300 65326 6302 65378
rect 6354 65326 6356 65378
rect 6300 64820 6356 65326
rect 6300 64596 6356 64764
rect 6300 64530 6356 64540
rect 6524 65266 6580 65660
rect 6636 65380 6692 66892
rect 6748 66836 6804 70140
rect 6860 67618 6916 67630
rect 6860 67566 6862 67618
rect 6914 67566 6916 67618
rect 6860 67508 6916 67566
rect 6860 67442 6916 67452
rect 6972 67058 7028 73500
rect 7196 73330 7252 73948
rect 7196 73278 7198 73330
rect 7250 73278 7252 73330
rect 7196 73266 7252 73278
rect 7084 73108 7140 73118
rect 7084 72770 7140 73052
rect 7084 72718 7086 72770
rect 7138 72718 7140 72770
rect 7084 72706 7140 72718
rect 7196 71764 7252 71774
rect 7196 71670 7252 71708
rect 7196 71540 7252 71550
rect 7084 70306 7140 70318
rect 7084 70254 7086 70306
rect 7138 70254 7140 70306
rect 7084 70196 7140 70254
rect 7196 70196 7252 71484
rect 7308 71202 7364 76412
rect 7532 75460 7588 76524
rect 7532 75394 7588 75404
rect 7532 74676 7588 74686
rect 7644 74676 7700 78204
rect 7980 75796 8036 75806
rect 8204 75796 8260 75806
rect 8036 75740 8148 75796
rect 7980 75730 8036 75740
rect 7756 75012 7812 75022
rect 7756 74918 7812 74956
rect 7644 74620 7812 74676
rect 7532 74582 7588 74620
rect 7644 74116 7700 74126
rect 7644 74022 7700 74060
rect 7756 74114 7812 74620
rect 7756 74062 7758 74114
rect 7810 74062 7812 74114
rect 7756 74050 7812 74062
rect 7868 74674 7924 74686
rect 7868 74622 7870 74674
rect 7922 74622 7924 74674
rect 7420 74002 7476 74014
rect 7420 73950 7422 74002
rect 7474 73950 7476 74002
rect 7420 73780 7476 73950
rect 7420 73714 7476 73724
rect 7644 73668 7700 73678
rect 7644 73554 7700 73612
rect 7644 73502 7646 73554
rect 7698 73502 7700 73554
rect 7644 73490 7700 73502
rect 7868 73556 7924 74622
rect 7980 74114 8036 74126
rect 7980 74062 7982 74114
rect 8034 74062 8036 74114
rect 7980 74004 8036 74062
rect 7980 73938 8036 73948
rect 8092 73948 8148 75740
rect 8204 75702 8260 75740
rect 8204 75348 8260 75358
rect 8204 74116 8260 75292
rect 8204 74050 8260 74060
rect 8092 73892 8260 73948
rect 7868 73490 7924 73500
rect 7868 73330 7924 73342
rect 7868 73278 7870 73330
rect 7922 73278 7924 73330
rect 7756 73218 7812 73230
rect 7756 73166 7758 73218
rect 7810 73166 7812 73218
rect 7420 73108 7476 73118
rect 7420 72770 7476 73052
rect 7420 72718 7422 72770
rect 7474 72718 7476 72770
rect 7420 72706 7476 72718
rect 7308 71150 7310 71202
rect 7362 71150 7364 71202
rect 7308 71138 7364 71150
rect 7420 71652 7476 71662
rect 7308 70980 7364 70990
rect 7308 70866 7364 70924
rect 7420 70978 7476 71596
rect 7420 70926 7422 70978
rect 7474 70926 7476 70978
rect 7420 70914 7476 70926
rect 7308 70814 7310 70866
rect 7362 70814 7364 70866
rect 7308 70532 7364 70814
rect 7308 70466 7364 70476
rect 7420 70644 7476 70654
rect 7084 70194 7252 70196
rect 7084 70142 7198 70194
rect 7250 70142 7252 70194
rect 7084 70140 7252 70142
rect 7196 70130 7252 70140
rect 7308 70084 7364 70094
rect 7308 69990 7364 70028
rect 7420 69636 7476 70588
rect 7532 70084 7588 70094
rect 7532 69990 7588 70028
rect 7196 69580 7476 69636
rect 7196 69522 7252 69580
rect 7196 69470 7198 69522
rect 7250 69470 7252 69522
rect 7196 69458 7252 69470
rect 7644 69410 7700 69422
rect 7644 69358 7646 69410
rect 7698 69358 7700 69410
rect 7196 68404 7252 68414
rect 7196 67954 7252 68348
rect 7196 67902 7198 67954
rect 7250 67902 7252 67954
rect 7196 67890 7252 67902
rect 6972 67006 6974 67058
rect 7026 67006 7028 67058
rect 6972 66994 7028 67006
rect 7084 67618 7140 67630
rect 7084 67566 7086 67618
rect 7138 67566 7140 67618
rect 6748 66780 7028 66836
rect 6748 66612 6804 66622
rect 6748 66386 6804 66556
rect 6748 66334 6750 66386
rect 6802 66334 6804 66386
rect 6748 66322 6804 66334
rect 6860 66164 6916 66174
rect 6860 66070 6916 66108
rect 6636 65314 6692 65324
rect 6748 65378 6804 65390
rect 6748 65326 6750 65378
rect 6802 65326 6804 65378
rect 6524 65214 6526 65266
rect 6578 65214 6580 65266
rect 6524 64594 6580 65214
rect 6748 65156 6804 65326
rect 6748 65090 6804 65100
rect 6524 64542 6526 64594
rect 6578 64542 6580 64594
rect 6524 64530 6580 64542
rect 6300 63922 6356 63934
rect 6300 63870 6302 63922
rect 6354 63870 6356 63922
rect 6300 63812 6356 63870
rect 6860 63924 6916 63934
rect 6860 63830 6916 63868
rect 6300 62916 6356 63756
rect 6860 63698 6916 63710
rect 6860 63646 6862 63698
rect 6914 63646 6916 63698
rect 6524 63362 6580 63374
rect 6524 63310 6526 63362
rect 6578 63310 6580 63362
rect 6524 63250 6580 63310
rect 6524 63198 6526 63250
rect 6578 63198 6580 63250
rect 6524 63186 6580 63198
rect 6636 63252 6692 63262
rect 6300 62850 6356 62860
rect 6412 62580 6468 62590
rect 6412 62486 6468 62524
rect 6188 62132 6468 62188
rect 6076 62066 6132 62076
rect 4956 61682 5124 61684
rect 4956 61630 4958 61682
rect 5010 61630 5124 61682
rect 4956 61628 5124 61630
rect 5852 61796 5908 61806
rect 5852 61682 5908 61740
rect 5852 61630 5854 61682
rect 5906 61630 5908 61682
rect 4956 61236 5012 61628
rect 5852 61618 5908 61630
rect 6300 61794 6356 61806
rect 6300 61742 6302 61794
rect 6354 61742 6356 61794
rect 6300 61682 6356 61742
rect 6300 61630 6302 61682
rect 6354 61630 6356 61682
rect 4956 61170 5012 61180
rect 5964 61572 6020 61582
rect 5292 61124 5348 61134
rect 4060 58548 4116 58558
rect 4172 58548 4228 58940
rect 4060 58546 4228 58548
rect 4060 58494 4062 58546
rect 4114 58494 4228 58546
rect 4060 58492 4228 58494
rect 4284 60674 4900 60676
rect 4284 60622 4510 60674
rect 4562 60622 4900 60674
rect 4284 60620 4900 60622
rect 4956 61012 5012 61022
rect 4060 58482 4116 58492
rect 3388 57810 3444 57820
rect 2940 57698 2996 57708
rect 2828 54450 2884 54460
rect 2716 49970 2772 49980
rect 4284 41860 4340 60620
rect 4508 60610 4564 60620
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4844 60226 4900 60238
rect 4844 60174 4846 60226
rect 4898 60174 4900 60226
rect 4844 60114 4900 60174
rect 4844 60062 4846 60114
rect 4898 60062 4900 60114
rect 4844 60050 4900 60062
rect 4396 60004 4452 60014
rect 4396 59780 4452 59948
rect 4396 59686 4452 59724
rect 4732 59892 4788 59902
rect 4732 59442 4788 59836
rect 4732 59390 4734 59442
rect 4786 59390 4788 59442
rect 4732 59378 4788 59390
rect 4844 59780 4900 59790
rect 4396 59108 4452 59118
rect 4396 59014 4452 59052
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4844 56868 4900 59724
rect 4956 59444 5012 60956
rect 4956 59378 5012 59388
rect 5292 59442 5348 61068
rect 5852 61124 5908 61134
rect 5852 61010 5908 61068
rect 5852 60958 5854 61010
rect 5906 60958 5908 61010
rect 5852 60946 5908 60958
rect 5516 60788 5572 60798
rect 5516 60694 5572 60732
rect 5852 59778 5908 59790
rect 5852 59726 5854 59778
rect 5906 59726 5908 59778
rect 5852 59556 5908 59726
rect 5852 59490 5908 59500
rect 5292 59390 5294 59442
rect 5346 59390 5348 59442
rect 5292 59378 5348 59390
rect 5964 59106 6020 61516
rect 6300 61348 6356 61630
rect 6300 61282 6356 61292
rect 6300 60788 6356 60798
rect 6300 60694 6356 60732
rect 6188 60116 6244 60126
rect 6188 59444 6244 60060
rect 6300 60004 6356 60014
rect 6300 59910 6356 59948
rect 6300 59444 6356 59454
rect 6188 59442 6356 59444
rect 6188 59390 6302 59442
rect 6354 59390 6356 59442
rect 6188 59388 6356 59390
rect 5964 59054 5966 59106
rect 6018 59054 6020 59106
rect 5852 58548 5908 58558
rect 5852 58454 5908 58492
rect 4844 56802 4900 56812
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5964 43652 6020 59054
rect 6076 58996 6132 59006
rect 6076 58902 6132 58940
rect 6300 58996 6356 59388
rect 6300 58930 6356 58940
rect 6300 58772 6356 58782
rect 6300 58546 6356 58716
rect 6300 58494 6302 58546
rect 6354 58494 6356 58546
rect 6300 58482 6356 58494
rect 6412 56308 6468 62132
rect 6636 61684 6692 63196
rect 6860 63252 6916 63646
rect 6860 63158 6916 63196
rect 6748 62242 6804 62254
rect 6748 62190 6750 62242
rect 6802 62190 6804 62242
rect 6748 61794 6804 62190
rect 6972 62188 7028 66780
rect 7084 66052 7140 67566
rect 7308 67620 7364 67630
rect 7308 67526 7364 67564
rect 7420 67172 7476 67182
rect 7420 67078 7476 67116
rect 7196 67058 7252 67070
rect 7196 67006 7198 67058
rect 7250 67006 7252 67058
rect 7196 66500 7252 67006
rect 7644 67058 7700 69358
rect 7644 67006 7646 67058
rect 7698 67006 7700 67058
rect 7308 66836 7364 66846
rect 7308 66742 7364 66780
rect 7196 66444 7364 66500
rect 7084 65986 7140 65996
rect 7196 66276 7252 66286
rect 7196 65716 7252 66220
rect 7308 66164 7364 66444
rect 7420 66164 7476 66174
rect 7308 66162 7476 66164
rect 7308 66110 7422 66162
rect 7474 66110 7476 66162
rect 7308 66108 7476 66110
rect 7420 65828 7476 66108
rect 7532 66052 7588 66062
rect 7532 65958 7588 65996
rect 7420 65772 7588 65828
rect 7196 65660 7476 65716
rect 7420 65658 7476 65660
rect 7420 65606 7422 65658
rect 7474 65606 7476 65658
rect 7420 65594 7476 65606
rect 7308 65546 7364 65558
rect 7308 65494 7310 65546
rect 7362 65494 7364 65546
rect 7084 65268 7140 65278
rect 7308 65268 7364 65494
rect 7084 65266 7364 65268
rect 7084 65214 7086 65266
rect 7138 65214 7364 65266
rect 7084 65212 7364 65214
rect 7084 65202 7140 65212
rect 7532 64708 7588 65772
rect 7644 65716 7700 67006
rect 7644 65650 7700 65660
rect 7420 64706 7588 64708
rect 7420 64654 7534 64706
rect 7586 64654 7588 64706
rect 7420 64652 7588 64654
rect 7196 64372 7252 64382
rect 7196 64146 7252 64316
rect 7196 64094 7198 64146
rect 7250 64094 7252 64146
rect 7196 63476 7252 64094
rect 7196 63410 7252 63420
rect 7308 63588 7364 63598
rect 7308 63364 7364 63532
rect 7308 63140 7364 63308
rect 7196 63084 7364 63140
rect 7196 62580 7252 63084
rect 7308 62916 7364 62926
rect 7308 62822 7364 62860
rect 7420 62580 7476 64652
rect 7532 64642 7588 64652
rect 7644 65490 7700 65502
rect 7644 65438 7646 65490
rect 7698 65438 7700 65490
rect 7644 64596 7700 65438
rect 7644 64530 7700 64540
rect 7756 64372 7812 73166
rect 7868 72324 7924 73278
rect 8204 72772 8260 73892
rect 8092 72716 8260 72772
rect 7980 72546 8036 72558
rect 7980 72494 7982 72546
rect 8034 72494 8036 72546
rect 7980 72436 8036 72494
rect 7980 72370 8036 72380
rect 7868 72258 7924 72268
rect 8092 72100 8148 72716
rect 8204 72548 8260 72558
rect 8204 72454 8260 72492
rect 7868 72044 8148 72100
rect 8204 72324 8260 72334
rect 7868 71540 7924 72044
rect 8092 71874 8148 71886
rect 8092 71822 8094 71874
rect 8146 71822 8148 71874
rect 7868 71474 7924 71484
rect 7980 71764 8036 71774
rect 7868 69412 7924 69422
rect 7868 69318 7924 69356
rect 7980 67954 8036 71708
rect 8092 70980 8148 71822
rect 8092 70914 8148 70924
rect 8092 70756 8148 70766
rect 8092 70662 8148 70700
rect 8204 70588 8260 72268
rect 8316 70756 8372 79324
rect 8876 79268 8932 79278
rect 8428 77812 8484 77822
rect 8428 76580 8484 77756
rect 8428 76514 8484 76524
rect 8876 76354 8932 79212
rect 8876 76302 8878 76354
rect 8930 76302 8932 76354
rect 8876 76290 8932 76302
rect 9100 77812 9156 77822
rect 8988 75684 9044 75694
rect 8988 75590 9044 75628
rect 8764 75460 8820 75470
rect 8652 75012 8708 75022
rect 8428 74898 8484 74910
rect 8428 74846 8430 74898
rect 8482 74846 8484 74898
rect 8428 74340 8484 74846
rect 8428 73332 8484 74284
rect 8540 74786 8596 74798
rect 8540 74734 8542 74786
rect 8594 74734 8596 74786
rect 8540 73668 8596 74734
rect 8652 74452 8708 74956
rect 8764 74900 8820 75404
rect 8764 74806 8820 74844
rect 8988 74900 9044 74910
rect 8988 74806 9044 74844
rect 8652 74396 8820 74452
rect 8652 74228 8708 74238
rect 8652 74114 8708 74172
rect 8652 74062 8654 74114
rect 8706 74062 8708 74114
rect 8652 74050 8708 74062
rect 8764 73668 8820 74396
rect 8876 74114 8932 74126
rect 8876 74062 8878 74114
rect 8930 74062 8932 74114
rect 8876 73892 8932 74062
rect 8876 73826 8932 73836
rect 8988 74002 9044 74014
rect 8988 73950 8990 74002
rect 9042 73950 9044 74002
rect 8988 73668 9044 73950
rect 8764 73612 8932 73668
rect 8540 73602 8596 73612
rect 8428 73276 8820 73332
rect 8540 73108 8596 73118
rect 8540 73014 8596 73052
rect 8652 73106 8708 73118
rect 8652 73054 8654 73106
rect 8706 73054 8708 73106
rect 8316 70690 8372 70700
rect 8428 72996 8484 73006
rect 8092 70532 8260 70588
rect 8092 69412 8148 70532
rect 8316 70420 8372 70430
rect 8316 70326 8372 70364
rect 8428 70308 8484 72940
rect 8652 72772 8708 73054
rect 8764 73108 8820 73276
rect 8876 73330 8932 73612
rect 8988 73602 9044 73612
rect 8988 73444 9044 73454
rect 9100 73444 9156 77756
rect 9660 77698 9716 77710
rect 9660 77646 9662 77698
rect 9714 77646 9716 77698
rect 9660 77252 9716 77646
rect 9548 75460 9604 75470
rect 8988 73442 9156 73444
rect 8988 73390 8990 73442
rect 9042 73390 9156 73442
rect 8988 73388 9156 73390
rect 9436 75458 9604 75460
rect 9436 75406 9550 75458
rect 9602 75406 9604 75458
rect 9436 75404 9604 75406
rect 9436 73892 9492 75404
rect 9548 75394 9604 75404
rect 9660 75236 9716 77196
rect 10220 77476 10276 77486
rect 9996 76916 10052 76926
rect 9996 76690 10052 76860
rect 9996 76638 9998 76690
rect 10050 76638 10052 76690
rect 9996 76626 10052 76638
rect 10108 75684 10164 75694
rect 10108 75590 10164 75628
rect 8988 73378 9044 73388
rect 8876 73278 8878 73330
rect 8930 73278 8932 73330
rect 8876 73266 8932 73278
rect 9324 73108 9380 73118
rect 8764 73052 9044 73108
rect 8652 72706 8708 72716
rect 8540 72324 8596 72334
rect 8540 72322 8708 72324
rect 8540 72270 8542 72322
rect 8594 72270 8708 72322
rect 8540 72268 8708 72270
rect 8540 72258 8596 72268
rect 8540 71652 8596 71662
rect 8540 71558 8596 71596
rect 8540 70420 8596 70430
rect 8540 70326 8596 70364
rect 8428 70242 8484 70252
rect 8204 70196 8260 70206
rect 8204 70102 8260 70140
rect 8428 70084 8484 70094
rect 8428 69990 8484 70028
rect 8204 69412 8260 69422
rect 8092 69356 8204 69412
rect 8204 69318 8260 69356
rect 8204 68516 8260 68526
rect 8204 68422 8260 68460
rect 7980 67902 7982 67954
rect 8034 67902 8036 67954
rect 7980 67890 8036 67902
rect 8428 67844 8484 67854
rect 8652 67844 8708 72268
rect 8876 71428 8932 71438
rect 8764 70194 8820 70206
rect 8764 70142 8766 70194
rect 8818 70142 8820 70194
rect 8764 70084 8820 70142
rect 8764 70018 8820 70028
rect 8876 69076 8932 71372
rect 8428 67842 8708 67844
rect 8428 67790 8430 67842
rect 8482 67790 8708 67842
rect 8428 67788 8708 67790
rect 8764 69020 8932 69076
rect 8428 67778 8484 67788
rect 7868 67730 7924 67742
rect 7868 67678 7870 67730
rect 7922 67678 7924 67730
rect 7868 66388 7924 67678
rect 8204 67730 8260 67742
rect 8764 67732 8820 69020
rect 8876 68852 8932 68862
rect 8876 68626 8932 68796
rect 8876 68574 8878 68626
rect 8930 68574 8932 68626
rect 8876 68562 8932 68574
rect 8204 67678 8206 67730
rect 8258 67678 8260 67730
rect 8204 66724 8260 67678
rect 8540 67676 8820 67732
rect 8876 68068 8932 68078
rect 8540 66946 8596 67676
rect 8876 67284 8932 68012
rect 8988 67730 9044 73052
rect 9100 72548 9156 72558
rect 9100 71428 9156 72492
rect 9100 71362 9156 71372
rect 9100 70420 9156 70430
rect 9100 69748 9156 70364
rect 9100 69298 9156 69692
rect 9100 69246 9102 69298
rect 9154 69246 9156 69298
rect 9100 69234 9156 69246
rect 9212 69636 9268 69646
rect 8988 67678 8990 67730
rect 9042 67678 9044 67730
rect 8988 67396 9044 67678
rect 8988 67330 9044 67340
rect 9100 67618 9156 67630
rect 9100 67566 9102 67618
rect 9154 67566 9156 67618
rect 8876 67190 8932 67228
rect 8764 67060 8820 67070
rect 8764 67058 8932 67060
rect 8764 67006 8766 67058
rect 8818 67006 8932 67058
rect 8764 67004 8932 67006
rect 8764 66994 8820 67004
rect 8540 66894 8542 66946
rect 8594 66894 8596 66946
rect 8204 66668 8484 66724
rect 8092 66500 8148 66510
rect 8092 66406 8148 66444
rect 8316 66500 8372 66510
rect 7868 66322 7924 66332
rect 8316 66162 8372 66444
rect 8316 66110 8318 66162
rect 8370 66110 8372 66162
rect 8316 66098 8372 66110
rect 8204 66052 8260 66062
rect 7980 66050 8260 66052
rect 7980 65998 8206 66050
rect 8258 65998 8260 66050
rect 7980 65996 8260 65998
rect 7868 64484 7924 64494
rect 7868 64390 7924 64428
rect 7196 62578 7364 62580
rect 7196 62526 7198 62578
rect 7250 62526 7364 62578
rect 7196 62524 7364 62526
rect 7196 62514 7252 62524
rect 6972 62132 7140 62188
rect 6748 61742 6750 61794
rect 6802 61742 6804 61794
rect 6748 61730 6804 61742
rect 6860 61908 6916 61918
rect 6636 61618 6692 61628
rect 6748 61572 6804 61582
rect 6860 61572 6916 61852
rect 6748 61570 6916 61572
rect 6748 61518 6750 61570
rect 6802 61518 6916 61570
rect 6748 61516 6916 61518
rect 6972 61796 7028 61806
rect 6748 61124 6804 61516
rect 6748 61058 6804 61068
rect 6860 61012 6916 61022
rect 6860 60918 6916 60956
rect 6636 59778 6692 59790
rect 6636 59726 6638 59778
rect 6690 59726 6692 59778
rect 6636 58994 6692 59726
rect 6860 59444 6916 59454
rect 6972 59444 7028 61740
rect 7084 60676 7140 62132
rect 7196 61684 7252 61694
rect 7196 61590 7252 61628
rect 7308 61236 7364 62524
rect 7420 62514 7476 62524
rect 7532 64316 7812 64372
rect 7308 61170 7364 61180
rect 7420 61794 7476 61806
rect 7420 61742 7422 61794
rect 7474 61742 7476 61794
rect 7196 60676 7252 60686
rect 7084 60620 7196 60676
rect 7196 60582 7252 60620
rect 7084 59780 7140 59790
rect 7084 59686 7140 59724
rect 6860 59442 7028 59444
rect 6860 59390 6862 59442
rect 6914 59390 7028 59442
rect 6860 59388 7028 59390
rect 7308 59444 7364 59454
rect 6860 59378 6916 59388
rect 7308 59350 7364 59388
rect 6636 58942 6638 58994
rect 6690 58942 6692 58994
rect 6636 58772 6692 58942
rect 6636 58706 6692 58716
rect 6412 56242 6468 56252
rect 6636 58212 6692 58222
rect 6748 58212 6804 58222
rect 6692 58210 6804 58212
rect 6692 58158 6750 58210
rect 6802 58158 6804 58210
rect 6692 58156 6804 58158
rect 6636 51940 6692 58156
rect 6748 58146 6804 58156
rect 7196 58210 7252 58222
rect 7196 58158 7198 58210
rect 7250 58158 7252 58210
rect 7196 58100 7252 58158
rect 7196 58034 7252 58044
rect 7308 57540 7364 57550
rect 7308 57446 7364 57484
rect 6636 51874 6692 51884
rect 7420 45220 7476 61742
rect 7532 61684 7588 64316
rect 7980 64036 8036 65996
rect 8204 65986 8260 65996
rect 8092 65716 8148 65726
rect 8092 64372 8148 65660
rect 8316 65716 8372 65726
rect 8316 65622 8372 65660
rect 8204 65604 8260 65614
rect 8204 65510 8260 65548
rect 8428 65492 8484 66668
rect 8316 65436 8484 65492
rect 8092 64306 8148 64316
rect 8204 64932 8260 64942
rect 8204 64146 8260 64876
rect 8204 64094 8206 64146
rect 8258 64094 8260 64146
rect 8204 64082 8260 64094
rect 7980 63980 8148 64036
rect 7644 63810 7700 63822
rect 7644 63758 7646 63810
rect 7698 63758 7700 63810
rect 7644 63588 7700 63758
rect 7980 63812 8036 63822
rect 7644 63522 7700 63532
rect 7756 63700 7812 63710
rect 7532 61618 7588 61628
rect 7644 62580 7700 62590
rect 7644 61348 7700 62524
rect 7756 62578 7812 63644
rect 7868 63140 7924 63150
rect 7868 63046 7924 63084
rect 7756 62526 7758 62578
rect 7810 62526 7812 62578
rect 7756 62514 7812 62526
rect 7980 62188 8036 63756
rect 8092 62580 8148 63980
rect 8092 62514 8148 62524
rect 8204 63476 8260 63486
rect 8204 63250 8260 63420
rect 8204 63198 8206 63250
rect 8258 63198 8260 63250
rect 8092 62354 8148 62366
rect 8092 62302 8094 62354
rect 8146 62302 8148 62354
rect 8092 62188 8148 62302
rect 7980 62132 8148 62188
rect 8204 62244 8260 63198
rect 8316 63252 8372 65436
rect 8540 65156 8596 66894
rect 8540 64932 8596 65100
rect 8540 64866 8596 64876
rect 8652 66612 8708 66622
rect 8316 63186 8372 63196
rect 8428 63812 8484 63822
rect 8428 62916 8484 63756
rect 8540 63700 8596 63710
rect 8540 63606 8596 63644
rect 8652 63362 8708 66556
rect 8876 66164 8932 67004
rect 8764 65492 8820 65502
rect 8764 65156 8820 65436
rect 8764 65090 8820 65100
rect 8764 64372 8820 64382
rect 8764 63922 8820 64316
rect 8764 63870 8766 63922
rect 8818 63870 8820 63922
rect 8764 63812 8820 63870
rect 8876 63924 8932 66108
rect 8988 66948 9044 66958
rect 8988 64708 9044 66892
rect 9100 66276 9156 67566
rect 9212 66386 9268 69580
rect 9324 68516 9380 73052
rect 9436 72660 9492 73836
rect 9436 72594 9492 72604
rect 9548 75180 9716 75236
rect 9548 70588 9604 75180
rect 9884 75012 9940 75022
rect 9660 74340 9716 74350
rect 9660 74246 9716 74284
rect 9772 74114 9828 74126
rect 9772 74062 9774 74114
rect 9826 74062 9828 74114
rect 9772 73948 9828 74062
rect 9884 74116 9940 74956
rect 9996 74674 10052 74686
rect 9996 74622 9998 74674
rect 10050 74622 10052 74674
rect 9996 74340 10052 74622
rect 9996 74274 10052 74284
rect 9996 74116 10052 74126
rect 9884 74114 10052 74116
rect 9884 74062 9998 74114
rect 10050 74062 10052 74114
rect 9884 74060 10052 74062
rect 9996 74050 10052 74060
rect 9436 70532 9604 70588
rect 9660 73892 9828 73948
rect 10108 74004 10164 74042
rect 10108 73938 10164 73948
rect 9660 70588 9716 73892
rect 9996 73780 10052 73790
rect 9996 72658 10052 73724
rect 10220 73780 10276 77420
rect 10444 76466 10500 76478
rect 10444 76414 10446 76466
rect 10498 76414 10500 76466
rect 10332 74676 10388 74686
rect 10332 74582 10388 74620
rect 10220 73714 10276 73724
rect 10444 73892 10500 76414
rect 10556 76466 10612 76478
rect 10556 76414 10558 76466
rect 10610 76414 10612 76466
rect 10556 75796 10612 76414
rect 10668 76466 10724 76478
rect 10668 76414 10670 76466
rect 10722 76414 10724 76466
rect 10668 76244 10724 76414
rect 10668 76178 10724 76188
rect 10892 76020 10948 79548
rect 11536 79200 11648 80000
rect 14364 79940 14420 79950
rect 10892 75954 10948 75964
rect 11452 77364 11508 77374
rect 10556 75730 10612 75740
rect 10668 75908 10724 75918
rect 10556 74788 10612 74798
rect 10556 74694 10612 74732
rect 10668 74114 10724 75852
rect 10780 75572 10836 75582
rect 10780 75570 10948 75572
rect 10780 75518 10782 75570
rect 10834 75518 10948 75570
rect 10780 75516 10948 75518
rect 10780 75506 10836 75516
rect 10668 74062 10670 74114
rect 10722 74062 10724 74114
rect 10668 74050 10724 74062
rect 10332 73668 10388 73678
rect 10220 73442 10276 73454
rect 10220 73390 10222 73442
rect 10274 73390 10276 73442
rect 10220 73332 10276 73390
rect 10220 73266 10276 73276
rect 10108 73220 10164 73230
rect 10108 73108 10164 73164
rect 10220 73108 10276 73118
rect 10108 73106 10276 73108
rect 10108 73054 10222 73106
rect 10274 73054 10276 73106
rect 10108 73052 10276 73054
rect 10220 73042 10276 73052
rect 9996 72606 9998 72658
rect 10050 72606 10052 72658
rect 9772 71988 9828 71998
rect 9772 71894 9828 71932
rect 9996 71764 10052 72606
rect 9660 70532 9940 70588
rect 9436 69636 9492 70532
rect 9436 69570 9492 69580
rect 9660 69860 9716 69870
rect 9660 69636 9716 69804
rect 9884 69860 9940 70532
rect 9996 70196 10052 71708
rect 10220 71540 10276 71550
rect 10220 71446 10276 71484
rect 10332 71092 10388 73612
rect 10444 72772 10500 73836
rect 10668 73780 10724 73790
rect 10668 73330 10724 73724
rect 10668 73278 10670 73330
rect 10722 73278 10724 73330
rect 10668 73220 10724 73278
rect 10668 73154 10724 73164
rect 10444 72706 10500 72716
rect 10892 72548 10948 75516
rect 11340 75460 11396 75470
rect 11340 75010 11396 75404
rect 11452 75348 11508 77308
rect 11564 77028 11620 79200
rect 12124 77588 12180 77598
rect 11788 77028 11844 77038
rect 11564 77026 11844 77028
rect 11564 76974 11790 77026
rect 11842 76974 11844 77026
rect 11564 76972 11844 76974
rect 11788 76962 11844 76972
rect 12012 76916 12068 76926
rect 11564 76692 11620 76702
rect 11564 76354 11620 76636
rect 11564 76302 11566 76354
rect 11618 76302 11620 76354
rect 11564 76132 11620 76302
rect 11564 76066 11620 76076
rect 11452 75292 11620 75348
rect 11340 74958 11342 75010
rect 11394 74958 11396 75010
rect 11340 74946 11396 74958
rect 11116 74900 11172 74910
rect 11116 74806 11172 74844
rect 11452 74898 11508 74910
rect 11452 74846 11454 74898
rect 11506 74846 11508 74898
rect 11228 74338 11284 74350
rect 11228 74286 11230 74338
rect 11282 74286 11284 74338
rect 11116 74228 11172 74238
rect 11004 74116 11060 74126
rect 11004 74022 11060 74060
rect 11116 74114 11172 74172
rect 11116 74062 11118 74114
rect 11170 74062 11172 74114
rect 11116 74050 11172 74062
rect 10668 72492 10948 72548
rect 10220 71036 10388 71092
rect 10556 72324 10612 72334
rect 9996 70130 10052 70140
rect 10108 70194 10164 70206
rect 10108 70142 10110 70194
rect 10162 70142 10164 70194
rect 9884 69794 9940 69804
rect 9548 69412 9604 69422
rect 9548 69318 9604 69356
rect 9324 68450 9380 68460
rect 9436 68964 9492 68974
rect 9324 68068 9380 68078
rect 9324 67842 9380 68012
rect 9324 67790 9326 67842
rect 9378 67790 9380 67842
rect 9324 67778 9380 67790
rect 9324 66612 9380 66622
rect 9324 66498 9380 66556
rect 9324 66446 9326 66498
rect 9378 66446 9380 66498
rect 9324 66434 9380 66446
rect 9212 66334 9214 66386
rect 9266 66334 9268 66386
rect 9212 66322 9268 66334
rect 9100 66210 9156 66220
rect 8988 64642 9044 64652
rect 9100 66050 9156 66062
rect 9100 65998 9102 66050
rect 9154 65998 9156 66050
rect 8988 64484 9044 64494
rect 8988 64390 9044 64428
rect 9100 64148 9156 65998
rect 9436 65940 9492 68908
rect 9660 68628 9716 69580
rect 9772 69300 9828 69310
rect 9772 68738 9828 69244
rect 9884 69188 9940 69198
rect 9884 68850 9940 69132
rect 9884 68798 9886 68850
rect 9938 68798 9940 68850
rect 9884 68786 9940 68798
rect 10108 68852 10164 70142
rect 10108 68786 10164 68796
rect 9772 68686 9774 68738
rect 9826 68686 9828 68738
rect 9772 68674 9828 68686
rect 9660 68562 9716 68572
rect 10108 68628 10164 68638
rect 10108 68292 10164 68572
rect 9996 68236 10164 68292
rect 9548 67730 9604 67742
rect 9548 67678 9550 67730
rect 9602 67678 9604 67730
rect 9548 67284 9604 67678
rect 9548 66836 9604 67228
rect 9548 66770 9604 66780
rect 9884 67508 9940 67518
rect 9100 64082 9156 64092
rect 9324 65884 9492 65940
rect 9660 66052 9716 66062
rect 8876 63868 9156 63924
rect 8764 63756 8932 63812
rect 8652 63310 8654 63362
rect 8706 63310 8708 63362
rect 8652 63298 8708 63310
rect 8764 63588 8820 63598
rect 8652 63140 8708 63150
rect 8764 63140 8820 63532
rect 8876 63364 8932 63756
rect 8876 63298 8932 63308
rect 8652 63138 8820 63140
rect 8652 63086 8654 63138
rect 8706 63086 8820 63138
rect 8652 63084 8820 63086
rect 8652 63074 8708 63084
rect 8428 62850 8484 62860
rect 8988 63028 9044 63038
rect 8540 62692 8596 62702
rect 8540 62580 8596 62636
rect 8204 62178 8260 62188
rect 8316 62578 8596 62580
rect 8316 62526 8542 62578
rect 8594 62526 8596 62578
rect 8316 62524 8596 62526
rect 8092 62020 8148 62132
rect 8316 62020 8372 62524
rect 8540 62514 8596 62524
rect 8988 62578 9044 62972
rect 8988 62526 8990 62578
rect 9042 62526 9044 62578
rect 8876 62244 8932 62254
rect 8092 61964 8372 62020
rect 8428 62130 8484 62142
rect 8428 62078 8430 62130
rect 8482 62078 8484 62130
rect 7756 61796 7812 61806
rect 7756 61684 7812 61740
rect 8428 61796 8484 62078
rect 8428 61730 8484 61740
rect 7756 61682 7924 61684
rect 7756 61630 7758 61682
rect 7810 61630 7924 61682
rect 7756 61628 7924 61630
rect 7756 61618 7812 61628
rect 7644 61282 7700 61292
rect 7756 60900 7812 60910
rect 7756 60806 7812 60844
rect 7756 60564 7812 60574
rect 7756 60228 7812 60508
rect 7868 60452 7924 61628
rect 8876 61682 8932 62188
rect 8876 61630 8878 61682
rect 8930 61630 8932 61682
rect 8876 61618 8932 61630
rect 8428 61348 8484 61358
rect 8316 61236 8372 61246
rect 7868 60386 7924 60396
rect 8092 60676 8148 60686
rect 7756 60114 7812 60172
rect 7756 60062 7758 60114
rect 7810 60062 7812 60114
rect 7756 60050 7812 60062
rect 8092 59780 8148 60620
rect 8204 60228 8260 60238
rect 8204 60114 8260 60172
rect 8204 60062 8206 60114
rect 8258 60062 8260 60114
rect 8204 60050 8260 60062
rect 7644 59556 7700 59566
rect 7644 59108 7700 59500
rect 8092 59332 8148 59724
rect 8092 59276 8260 59332
rect 7980 59220 8036 59230
rect 8036 59164 8148 59220
rect 7644 59106 7812 59108
rect 7644 59054 7646 59106
rect 7698 59054 7812 59106
rect 7644 59052 7812 59054
rect 7644 59042 7700 59052
rect 7644 58212 7700 58222
rect 7644 58118 7700 58156
rect 7756 53732 7812 59052
rect 7868 57876 7924 57886
rect 7868 57782 7924 57820
rect 7980 56532 8036 59164
rect 8092 59106 8148 59164
rect 8092 59054 8094 59106
rect 8146 59054 8148 59106
rect 8092 59042 8148 59054
rect 7980 56466 8036 56476
rect 8092 58210 8148 58222
rect 8092 58158 8094 58210
rect 8146 58158 8148 58210
rect 8092 57316 8148 58158
rect 8092 55300 8148 57260
rect 8204 57092 8260 59276
rect 8316 57874 8372 61180
rect 8428 60564 8484 61292
rect 8652 61124 8708 61134
rect 8652 61010 8708 61068
rect 8652 60958 8654 61010
rect 8706 60958 8708 61010
rect 8652 60788 8708 60958
rect 8988 61012 9044 62526
rect 8988 60946 9044 60956
rect 8652 60722 8708 60732
rect 8428 60498 8484 60508
rect 8988 60674 9044 60686
rect 8988 60622 8990 60674
rect 9042 60622 9044 60674
rect 8988 60564 9044 60622
rect 8988 60498 9044 60508
rect 8652 60228 8708 60238
rect 8652 60114 8708 60172
rect 9100 60228 9156 63868
rect 9212 63700 9268 63710
rect 9212 63140 9268 63644
rect 9324 63476 9380 65884
rect 9436 65380 9492 65390
rect 9436 64706 9492 65324
rect 9436 64654 9438 64706
rect 9490 64654 9492 64706
rect 9436 64642 9492 64654
rect 9660 64594 9716 65996
rect 9660 64542 9662 64594
rect 9714 64542 9716 64594
rect 9660 64530 9716 64542
rect 9772 64594 9828 64606
rect 9772 64542 9774 64594
rect 9826 64542 9828 64594
rect 9548 64482 9604 64494
rect 9548 64430 9550 64482
rect 9602 64430 9604 64482
rect 9548 63700 9604 64430
rect 9772 64372 9828 64542
rect 9884 64596 9940 67452
rect 9996 66050 10052 68236
rect 10108 68068 10164 68078
rect 10108 67842 10164 68012
rect 10220 67954 10276 71036
rect 10332 70866 10388 70878
rect 10332 70814 10334 70866
rect 10386 70814 10388 70866
rect 10332 70644 10388 70814
rect 10332 70578 10388 70588
rect 10444 70308 10500 70318
rect 10332 69410 10388 69422
rect 10332 69358 10334 69410
rect 10386 69358 10388 69410
rect 10332 68404 10388 69358
rect 10444 68964 10500 70252
rect 10556 70084 10612 72268
rect 10668 72100 10724 72492
rect 11004 72436 11060 72446
rect 11004 72342 11060 72380
rect 11116 72434 11172 72446
rect 11116 72382 11118 72434
rect 11170 72382 11172 72434
rect 10780 72324 10836 72334
rect 11116 72324 11172 72382
rect 10780 72322 10948 72324
rect 10780 72270 10782 72322
rect 10834 72270 10948 72322
rect 10780 72268 10948 72270
rect 10780 72258 10836 72268
rect 10668 72034 10724 72044
rect 10892 72100 10948 72268
rect 11116 72258 11172 72268
rect 10892 72034 10948 72044
rect 10668 71764 10724 71774
rect 10668 71670 10724 71708
rect 10780 71762 10836 71774
rect 10780 71710 10782 71762
rect 10834 71710 10836 71762
rect 10780 71316 10836 71710
rect 10780 71250 10836 71260
rect 10892 71762 10948 71774
rect 10892 71710 10894 71762
rect 10946 71710 10948 71762
rect 10892 71092 10948 71710
rect 10892 71026 10948 71036
rect 11004 70978 11060 70990
rect 11004 70926 11006 70978
rect 11058 70926 11060 70978
rect 10780 70084 10836 70094
rect 10556 70082 10836 70084
rect 10556 70030 10782 70082
rect 10834 70030 10836 70082
rect 10556 70028 10836 70030
rect 10668 69748 10724 69758
rect 10444 68908 10612 68964
rect 10444 68628 10500 68638
rect 10444 68534 10500 68572
rect 10332 68338 10388 68348
rect 10220 67902 10222 67954
rect 10274 67902 10276 67954
rect 10220 67890 10276 67902
rect 10332 68180 10388 68190
rect 10108 67790 10110 67842
rect 10162 67790 10164 67842
rect 10108 67778 10164 67790
rect 10332 67842 10388 68124
rect 10332 67790 10334 67842
rect 10386 67790 10388 67842
rect 10332 67778 10388 67790
rect 10556 67730 10612 68908
rect 10668 68628 10724 69692
rect 10780 68964 10836 70028
rect 10892 69188 10948 69198
rect 10892 69094 10948 69132
rect 10780 68898 10836 68908
rect 11004 68852 11060 70926
rect 11004 68786 11060 68796
rect 11116 70756 11172 70766
rect 10668 68562 10724 68572
rect 10892 68628 10948 68638
rect 10556 67678 10558 67730
rect 10610 67678 10612 67730
rect 10556 67284 10612 67678
rect 10556 67218 10612 67228
rect 10668 68402 10724 68414
rect 10892 68404 10948 68572
rect 10668 68350 10670 68402
rect 10722 68350 10724 68402
rect 10108 67170 10164 67182
rect 10108 67118 10110 67170
rect 10162 67118 10164 67170
rect 10108 66948 10164 67118
rect 10668 67172 10724 68350
rect 10668 67106 10724 67116
rect 10780 68402 10948 68404
rect 10780 68350 10894 68402
rect 10946 68350 10948 68402
rect 10780 68348 10948 68350
rect 10108 66882 10164 66892
rect 10332 67058 10388 67070
rect 10332 67006 10334 67058
rect 10386 67006 10388 67058
rect 9996 65998 9998 66050
rect 10050 65998 10052 66050
rect 9996 65986 10052 65998
rect 10220 65604 10276 65614
rect 10332 65604 10388 67006
rect 10556 67058 10612 67070
rect 10556 67006 10558 67058
rect 10610 67006 10612 67058
rect 10220 65602 10388 65604
rect 10220 65550 10222 65602
rect 10274 65550 10388 65602
rect 10220 65548 10388 65550
rect 10444 66946 10500 66958
rect 10444 66894 10446 66946
rect 10498 66894 10500 66946
rect 10444 65604 10500 66894
rect 10556 66948 10612 67006
rect 10556 66882 10612 66892
rect 10556 66276 10612 66286
rect 10556 66182 10612 66220
rect 10220 65380 10276 65548
rect 10444 65538 10500 65548
rect 10556 65940 10612 65950
rect 10108 65266 10164 65278
rect 10108 65214 10110 65266
rect 10162 65214 10164 65266
rect 10108 65044 10164 65214
rect 10108 64978 10164 64988
rect 9996 64596 10052 64606
rect 9884 64594 10052 64596
rect 9884 64542 9998 64594
rect 10050 64542 10052 64594
rect 9884 64540 10052 64542
rect 9996 64530 10052 64540
rect 10108 64596 10164 64606
rect 10108 64372 10164 64540
rect 9772 64316 10164 64372
rect 9548 63634 9604 63644
rect 9996 63924 10052 63934
rect 9996 63476 10052 63868
rect 9324 63420 9716 63476
rect 9212 63008 9268 63084
rect 9324 62916 9380 62926
rect 9100 60162 9156 60172
rect 9212 62244 9268 62254
rect 8652 60062 8654 60114
rect 8706 60062 8708 60114
rect 8652 60050 8708 60062
rect 8988 60116 9044 60126
rect 8652 59556 8708 59566
rect 8652 59442 8708 59500
rect 8652 59390 8654 59442
rect 8706 59390 8708 59442
rect 8652 59378 8708 59390
rect 8988 59332 9044 60060
rect 9100 59444 9156 59454
rect 9100 59350 9156 59388
rect 8988 59266 9044 59276
rect 9212 58828 9268 62188
rect 9324 61682 9380 62860
rect 9548 62914 9604 62926
rect 9548 62862 9550 62914
rect 9602 62862 9604 62914
rect 9548 62020 9604 62862
rect 9548 61954 9604 61964
rect 9324 61630 9326 61682
rect 9378 61630 9380 61682
rect 9324 61618 9380 61630
rect 9436 60116 9492 60126
rect 9436 60022 9492 60060
rect 9660 59444 9716 63420
rect 9996 63410 10052 63420
rect 10220 63364 10276 65324
rect 10332 65268 10388 65278
rect 10332 65044 10388 65212
rect 10332 64978 10388 64988
rect 10444 65266 10500 65278
rect 10444 65214 10446 65266
rect 10498 65214 10500 65266
rect 10444 64820 10500 65214
rect 10444 64754 10500 64764
rect 10332 63812 10388 63822
rect 10332 63718 10388 63756
rect 10332 63364 10388 63374
rect 10220 63362 10388 63364
rect 10220 63310 10334 63362
rect 10386 63310 10388 63362
rect 10220 63308 10388 63310
rect 9996 63252 10052 63262
rect 9996 63158 10052 63196
rect 10108 63140 10164 63150
rect 9996 62244 10052 62254
rect 10108 62244 10164 63084
rect 10220 62692 10276 63308
rect 10332 63298 10388 63308
rect 10556 63250 10612 65884
rect 10556 63198 10558 63250
rect 10610 63198 10612 63250
rect 10556 63028 10612 63198
rect 10780 63140 10836 68348
rect 10892 68338 10948 68348
rect 11004 68404 11060 68414
rect 11004 68310 11060 68348
rect 11116 68180 11172 70700
rect 10780 63074 10836 63084
rect 10892 68124 11172 68180
rect 10892 66500 10948 68124
rect 11228 67956 11284 74286
rect 11452 74340 11508 74846
rect 11452 74274 11508 74284
rect 11340 74114 11396 74126
rect 11340 74062 11342 74114
rect 11394 74062 11396 74114
rect 11340 74004 11396 74062
rect 11340 73668 11396 73948
rect 11340 73602 11396 73612
rect 11340 73330 11396 73342
rect 11340 73278 11342 73330
rect 11394 73278 11396 73330
rect 11340 72548 11396 73278
rect 11340 72482 11396 72492
rect 11452 73332 11508 73342
rect 10892 64482 10948 66444
rect 11116 67900 11284 67956
rect 11340 71764 11396 71774
rect 11340 69300 11396 71708
rect 11452 70308 11508 73276
rect 11564 72324 11620 75292
rect 11900 74674 11956 74686
rect 11900 74622 11902 74674
rect 11954 74622 11956 74674
rect 11788 74452 11844 74462
rect 11788 74338 11844 74396
rect 11788 74286 11790 74338
rect 11842 74286 11844 74338
rect 11788 74004 11844 74286
rect 11788 73938 11844 73948
rect 11900 73892 11956 74622
rect 12012 74340 12068 76860
rect 12124 76692 12180 77532
rect 12124 75908 12180 76636
rect 12124 75842 12180 75852
rect 12236 77476 12292 77486
rect 12236 74452 12292 77420
rect 13804 77364 13860 77374
rect 12348 77026 12404 77038
rect 12348 76974 12350 77026
rect 12402 76974 12404 77026
rect 12348 76580 12404 76974
rect 12348 76578 12516 76580
rect 12348 76526 12350 76578
rect 12402 76526 12516 76578
rect 12348 76524 12516 76526
rect 12348 76514 12404 76524
rect 12348 75908 12404 75918
rect 12348 75122 12404 75852
rect 12348 75070 12350 75122
rect 12402 75070 12404 75122
rect 12348 75058 12404 75070
rect 12460 74676 12516 76524
rect 13580 76356 13636 76366
rect 13468 75908 13524 75918
rect 12908 75796 12964 75806
rect 12908 75702 12964 75740
rect 13132 75124 13188 75134
rect 13020 75012 13076 75022
rect 13020 74918 13076 74956
rect 13132 75010 13188 75068
rect 13132 74958 13134 75010
rect 13186 74958 13188 75010
rect 13132 74946 13188 74958
rect 12460 74610 12516 74620
rect 12572 74898 12628 74910
rect 12572 74846 12574 74898
rect 12626 74846 12628 74898
rect 12236 74396 12516 74452
rect 12012 74284 12404 74340
rect 12012 74116 12068 74126
rect 12012 74022 12068 74060
rect 11788 73220 11844 73230
rect 11676 72884 11732 72894
rect 11676 72658 11732 72828
rect 11676 72606 11678 72658
rect 11730 72606 11732 72658
rect 11676 72594 11732 72606
rect 11564 72258 11620 72268
rect 11452 70242 11508 70252
rect 11676 71652 11732 71662
rect 11564 69300 11620 69310
rect 11340 69298 11620 69300
rect 11340 69246 11566 69298
rect 11618 69246 11620 69298
rect 11340 69244 11620 69246
rect 11116 66388 11172 67900
rect 11228 67732 11284 67742
rect 11228 67638 11284 67676
rect 11340 66948 11396 69244
rect 11564 69234 11620 69244
rect 11676 69300 11732 71596
rect 11788 70756 11844 73164
rect 11900 72996 11956 73836
rect 11900 72930 11956 72940
rect 12124 74004 12180 74014
rect 12012 72658 12068 72670
rect 12012 72606 12014 72658
rect 12066 72606 12068 72658
rect 11900 71876 11956 71886
rect 11900 71090 11956 71820
rect 11900 71038 11902 71090
rect 11954 71038 11956 71090
rect 11900 71026 11956 71038
rect 11788 70690 11844 70700
rect 11676 69168 11732 69244
rect 11900 69186 11956 69198
rect 11900 69134 11902 69186
rect 11954 69134 11956 69186
rect 11564 68852 11620 68862
rect 11564 68516 11620 68796
rect 11788 68516 11844 68526
rect 11564 68514 11844 68516
rect 11564 68462 11790 68514
rect 11842 68462 11844 68514
rect 11564 68460 11844 68462
rect 11340 66882 11396 66892
rect 11452 68292 11508 68302
rect 11452 67842 11508 68236
rect 11452 67790 11454 67842
rect 11506 67790 11508 67842
rect 11452 66724 11508 67790
rect 11564 67060 11620 68460
rect 11788 68450 11844 68460
rect 11676 68292 11732 68302
rect 11676 67954 11732 68236
rect 11900 68292 11956 69134
rect 11900 68226 11956 68236
rect 11676 67902 11678 67954
rect 11730 67902 11732 67954
rect 11676 67890 11732 67902
rect 11788 67732 11844 67742
rect 11788 67638 11844 67676
rect 11564 67058 11732 67060
rect 11564 67006 11566 67058
rect 11618 67006 11732 67058
rect 11564 67004 11732 67006
rect 11564 66994 11620 67004
rect 11452 66658 11508 66668
rect 11116 66322 11172 66332
rect 11564 66164 11620 66174
rect 11564 66070 11620 66108
rect 11228 65492 11284 65502
rect 10892 64430 10894 64482
rect 10946 64430 10948 64482
rect 10556 62962 10612 62972
rect 10220 62626 10276 62636
rect 10780 62580 10836 62590
rect 10780 62486 10836 62524
rect 10668 62468 10724 62478
rect 10052 62188 10164 62244
rect 10556 62354 10612 62366
rect 10556 62302 10558 62354
rect 10610 62302 10612 62354
rect 9996 62150 10052 62188
rect 9772 62132 9828 62142
rect 9772 60788 9828 62076
rect 10556 61908 10612 62302
rect 10668 62244 10724 62412
rect 10668 62178 10724 62188
rect 10892 62188 10948 64430
rect 11116 65378 11172 65390
rect 11116 65326 11118 65378
rect 11170 65326 11172 65378
rect 11116 62804 11172 65326
rect 11228 63924 11284 65436
rect 11564 64482 11620 64494
rect 11564 64430 11566 64482
rect 11618 64430 11620 64482
rect 11452 64260 11508 64270
rect 11452 64146 11508 64204
rect 11452 64094 11454 64146
rect 11506 64094 11508 64146
rect 11452 64082 11508 64094
rect 11228 63858 11284 63868
rect 11340 63812 11396 63822
rect 11340 63364 11396 63756
rect 11340 63138 11396 63308
rect 11564 63364 11620 64430
rect 11564 63298 11620 63308
rect 11340 63086 11342 63138
rect 11394 63086 11396 63138
rect 11340 63074 11396 63086
rect 11676 63028 11732 67004
rect 11900 66386 11956 66398
rect 11900 66334 11902 66386
rect 11954 66334 11956 66386
rect 11900 65380 11956 66334
rect 11900 65314 11956 65324
rect 12012 65156 12068 72606
rect 12124 69524 12180 73948
rect 12236 72548 12292 72558
rect 12236 72454 12292 72492
rect 12348 69972 12404 74284
rect 12460 72324 12516 74396
rect 12572 73108 12628 74846
rect 13356 74788 13412 74798
rect 13132 74676 13188 74686
rect 12684 74172 13076 74228
rect 12684 74002 12740 74172
rect 12684 73950 12686 74002
rect 12738 73950 12740 74002
rect 12684 73938 12740 73950
rect 12796 74004 12852 74042
rect 12796 73938 12852 73948
rect 12908 74002 12964 74014
rect 12908 73950 12910 74002
rect 12962 73950 12964 74002
rect 12796 73220 12852 73230
rect 12796 73126 12852 73164
rect 12572 73042 12628 73052
rect 12908 72436 12964 73950
rect 13020 73332 13076 74172
rect 13020 73200 13076 73276
rect 12908 72370 12964 72380
rect 12460 72268 12852 72324
rect 12684 71316 12740 71326
rect 12572 70980 12628 70990
rect 12460 70754 12516 70766
rect 12460 70702 12462 70754
rect 12514 70702 12516 70754
rect 12460 70644 12516 70702
rect 12460 70578 12516 70588
rect 12572 70644 12628 70924
rect 12684 70978 12740 71260
rect 12796 71090 12852 72268
rect 12796 71038 12798 71090
rect 12850 71038 12852 71090
rect 12796 71026 12852 71038
rect 12684 70926 12686 70978
rect 12738 70926 12740 70978
rect 12684 70914 12740 70926
rect 13020 70980 13076 70990
rect 12908 70756 12964 70766
rect 12908 70662 12964 70700
rect 12684 70644 12740 70654
rect 12572 70588 12684 70644
rect 12572 70196 12628 70588
rect 12684 70578 12740 70588
rect 12572 70140 12964 70196
rect 12908 70082 12964 70140
rect 12908 70030 12910 70082
rect 12962 70030 12964 70082
rect 12908 70018 12964 70030
rect 12348 69916 12852 69972
rect 12684 69524 12740 69534
rect 12180 69468 12292 69524
rect 12124 69392 12180 69468
rect 11788 65100 12068 65156
rect 12124 69188 12180 69198
rect 12236 69188 12292 69468
rect 12460 69412 12516 69422
rect 12684 69412 12740 69468
rect 12460 69410 12740 69412
rect 12460 69358 12462 69410
rect 12514 69358 12740 69410
rect 12460 69356 12740 69358
rect 12460 69346 12516 69356
rect 12348 69188 12404 69198
rect 12236 69186 12404 69188
rect 12236 69134 12350 69186
rect 12402 69134 12404 69186
rect 12236 69132 12404 69134
rect 11788 64148 11844 65100
rect 11900 64932 11956 64942
rect 12124 64932 12180 69132
rect 12348 69122 12404 69132
rect 12572 69186 12628 69198
rect 12572 69134 12574 69186
rect 12626 69134 12628 69186
rect 12572 69076 12628 69134
rect 12572 68964 12628 69020
rect 12348 68908 12628 68964
rect 12236 66948 12292 66958
rect 12236 66854 12292 66892
rect 11900 64930 12180 64932
rect 11900 64878 11902 64930
rect 11954 64878 12180 64930
rect 11900 64876 12180 64878
rect 11900 64866 11956 64876
rect 12124 64708 12180 64718
rect 12124 64594 12180 64652
rect 12124 64542 12126 64594
rect 12178 64542 12180 64594
rect 12124 64530 12180 64542
rect 12348 64596 12404 68908
rect 12796 68852 12852 69916
rect 13020 69410 13076 70924
rect 13020 69358 13022 69410
rect 13074 69358 13076 69410
rect 13020 69346 13076 69358
rect 12460 68796 12852 68852
rect 12460 68066 12516 68796
rect 12684 68628 12740 68638
rect 12908 68628 12964 68638
rect 12740 68572 12852 68628
rect 12684 68562 12740 68572
rect 12460 68014 12462 68066
rect 12514 68014 12516 68066
rect 12460 68002 12516 68014
rect 12796 68066 12852 68572
rect 12796 68014 12798 68066
rect 12850 68014 12852 68066
rect 12796 68002 12852 68014
rect 12908 68066 12964 68572
rect 12908 68014 12910 68066
rect 12962 68014 12964 68066
rect 12908 68002 12964 68014
rect 12684 67956 12740 67966
rect 12572 67842 12628 67854
rect 12572 67790 12574 67842
rect 12626 67790 12628 67842
rect 12572 67396 12628 67790
rect 12572 67330 12628 67340
rect 12684 67060 12740 67900
rect 12684 66274 12740 67004
rect 12684 66222 12686 66274
rect 12738 66222 12740 66274
rect 12684 66210 12740 66222
rect 12796 67284 12852 67294
rect 12796 66052 12852 67228
rect 12684 65996 12796 66052
rect 12460 65716 12516 65726
rect 12460 65602 12516 65660
rect 12460 65550 12462 65602
rect 12514 65550 12516 65602
rect 12460 65538 12516 65550
rect 12348 64530 12404 64540
rect 12572 64594 12628 64606
rect 12572 64542 12574 64594
rect 12626 64542 12628 64594
rect 12572 64484 12628 64542
rect 12460 64428 12572 64484
rect 12124 64148 12180 64158
rect 11788 64146 12180 64148
rect 11788 64094 12126 64146
rect 12178 64094 12180 64146
rect 11788 64092 12180 64094
rect 12124 64082 12180 64092
rect 12348 64036 12404 64046
rect 12460 64036 12516 64428
rect 12572 64418 12628 64428
rect 12348 64034 12516 64036
rect 12348 63982 12350 64034
rect 12402 63982 12516 64034
rect 12348 63980 12516 63982
rect 11900 63924 11956 63934
rect 11116 62738 11172 62748
rect 11452 62972 11732 63028
rect 11788 63588 11844 63598
rect 11228 62356 11284 62366
rect 11228 62262 11284 62300
rect 10780 62132 10836 62142
rect 10892 62132 11396 62188
rect 10780 61908 10836 62076
rect 10780 61852 10948 61908
rect 10556 61842 10612 61852
rect 9884 61684 9940 61694
rect 9884 61590 9940 61628
rect 10780 61684 10836 61694
rect 10780 61590 10836 61628
rect 10892 61682 10948 61852
rect 10892 61630 10894 61682
rect 10946 61630 10948 61682
rect 10892 61618 10948 61630
rect 10220 61572 10276 61582
rect 10220 61478 10276 61516
rect 11116 61572 11172 61582
rect 11116 61478 11172 61516
rect 9772 60722 9828 60732
rect 9884 61460 9940 61470
rect 9884 60564 9940 61404
rect 10108 61124 10164 61134
rect 10108 61010 10164 61068
rect 10108 60958 10110 61010
rect 10162 60958 10164 61010
rect 10108 60946 10164 60958
rect 10220 61012 10276 61022
rect 10220 60918 10276 60956
rect 10780 61012 10836 61022
rect 10780 60918 10836 60956
rect 11116 61012 11172 61022
rect 9996 60564 10052 60574
rect 9940 60562 10052 60564
rect 9940 60510 9998 60562
rect 10050 60510 10052 60562
rect 9940 60508 10052 60510
rect 9884 60432 9940 60508
rect 9996 60498 10052 60508
rect 10668 60564 10724 60574
rect 10668 60114 10724 60508
rect 10668 60062 10670 60114
rect 10722 60062 10724 60114
rect 10668 60050 10724 60062
rect 9996 59892 10052 59902
rect 9884 59836 9996 59892
rect 9772 59444 9828 59454
rect 9660 59442 9828 59444
rect 9660 59390 9774 59442
rect 9826 59390 9828 59442
rect 9660 59388 9828 59390
rect 9772 59378 9828 59388
rect 9772 59220 9828 59230
rect 9212 58772 9380 58828
rect 9324 58546 9380 58716
rect 9324 58494 9326 58546
rect 9378 58494 9380 58546
rect 9324 58482 9380 58494
rect 9772 58546 9828 59164
rect 9772 58494 9774 58546
rect 9826 58494 9828 58546
rect 9772 58482 9828 58494
rect 8316 57822 8318 57874
rect 8370 57822 8372 57874
rect 8316 57810 8372 57822
rect 8764 58210 8820 58222
rect 8764 58158 8766 58210
rect 8818 58158 8820 58210
rect 8764 57764 8820 58158
rect 8988 57876 9044 57886
rect 8988 57782 9044 57820
rect 9772 57876 9828 57886
rect 9884 57876 9940 59836
rect 9996 59798 10052 59836
rect 10556 59668 10612 59678
rect 10444 59220 10500 59230
rect 10220 59108 10276 59118
rect 10444 59108 10500 59164
rect 10220 58546 10276 59052
rect 10220 58494 10222 58546
rect 10274 58494 10276 58546
rect 10220 58482 10276 58494
rect 10332 59106 10500 59108
rect 10332 59054 10446 59106
rect 10498 59054 10500 59106
rect 10332 59052 10500 59054
rect 9772 57874 9940 57876
rect 9772 57822 9774 57874
rect 9826 57822 9940 57874
rect 9772 57820 9940 57822
rect 9772 57810 9828 57820
rect 8764 57698 8820 57708
rect 10220 57540 10276 57550
rect 8204 57026 8260 57036
rect 9996 57092 10052 57102
rect 9324 56980 9380 56990
rect 9324 56756 9380 56924
rect 9772 56980 9828 56990
rect 9772 56886 9828 56924
rect 9324 56690 9380 56700
rect 8092 55234 8148 55244
rect 7756 53666 7812 53676
rect 8316 53732 8372 53742
rect 7420 45154 7476 45164
rect 8204 45220 8260 45230
rect 5964 43586 6020 43596
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4284 41794 4340 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 8204 5908 8260 45164
rect 8316 6020 8372 53676
rect 8316 5954 8372 5964
rect 9996 48356 10052 57036
rect 10220 56978 10276 57484
rect 10220 56926 10222 56978
rect 10274 56926 10276 56978
rect 10220 56914 10276 56926
rect 10332 52052 10388 59052
rect 10444 59042 10500 59052
rect 10444 57876 10500 57886
rect 10556 57876 10612 59612
rect 10780 59108 10836 59118
rect 10780 59014 10836 59052
rect 10668 58436 10724 58446
rect 10668 58342 10724 58380
rect 10444 57874 10612 57876
rect 10444 57822 10446 57874
rect 10498 57822 10612 57874
rect 10444 57820 10612 57822
rect 11116 57876 11172 60956
rect 11228 60228 11284 60238
rect 11228 60114 11284 60172
rect 11228 60062 11230 60114
rect 11282 60062 11284 60114
rect 11228 60050 11284 60062
rect 11228 59444 11284 59454
rect 11228 59350 11284 59388
rect 11340 59108 11396 62132
rect 11452 60900 11508 62972
rect 11564 62804 11620 62814
rect 11564 61682 11620 62748
rect 11676 62468 11732 62478
rect 11788 62468 11844 63532
rect 11900 63028 11956 63868
rect 12012 63922 12068 63934
rect 12012 63870 12014 63922
rect 12066 63870 12068 63922
rect 12012 63588 12068 63870
rect 12348 63812 12404 63980
rect 12348 63746 12404 63756
rect 12012 63250 12068 63532
rect 12012 63198 12014 63250
rect 12066 63198 12068 63250
rect 12012 63186 12068 63198
rect 12236 63140 12292 63150
rect 12292 63084 12404 63140
rect 12236 63046 12292 63084
rect 11900 62972 12068 63028
rect 11676 62466 11844 62468
rect 11676 62414 11678 62466
rect 11730 62414 11844 62466
rect 11676 62412 11844 62414
rect 11676 62402 11732 62412
rect 11788 62188 11844 62412
rect 11900 62692 11956 62702
rect 11900 62354 11956 62636
rect 11900 62302 11902 62354
rect 11954 62302 11956 62354
rect 11900 62290 11956 62302
rect 11788 62132 11956 62188
rect 11564 61630 11566 61682
rect 11618 61630 11620 61682
rect 11564 61618 11620 61630
rect 11900 61460 11956 62132
rect 12012 61572 12068 62972
rect 12012 61506 12068 61516
rect 12124 62916 12180 62926
rect 12124 62580 12180 62860
rect 12236 62580 12292 62590
rect 12124 62578 12292 62580
rect 12124 62526 12238 62578
rect 12290 62526 12292 62578
rect 12124 62524 12292 62526
rect 11452 60844 11620 60900
rect 11228 58548 11284 58558
rect 11340 58548 11396 59052
rect 11452 60674 11508 60686
rect 11452 60622 11454 60674
rect 11506 60622 11508 60674
rect 11452 60452 11508 60622
rect 11452 59444 11508 60396
rect 11452 58996 11508 59388
rect 11452 58930 11508 58940
rect 11564 60116 11620 60844
rect 11900 60674 11956 61404
rect 11900 60622 11902 60674
rect 11954 60622 11956 60674
rect 11900 60564 11956 60622
rect 11900 60498 11956 60508
rect 12012 61348 12068 61358
rect 11228 58546 11396 58548
rect 11228 58494 11230 58546
rect 11282 58494 11396 58546
rect 11228 58492 11396 58494
rect 11564 58548 11620 60060
rect 11676 60228 11732 60238
rect 11676 60002 11732 60172
rect 11676 59950 11678 60002
rect 11730 59950 11732 60002
rect 11676 59938 11732 59950
rect 12012 60228 12068 61292
rect 12124 60340 12180 62524
rect 12236 62514 12292 62524
rect 12348 61796 12404 63084
rect 12460 62130 12516 63980
rect 12460 62078 12462 62130
rect 12514 62078 12516 62130
rect 12460 62066 12516 62078
rect 12572 63924 12628 63934
rect 12348 61740 12516 61796
rect 12348 61572 12404 61582
rect 12460 61572 12516 61740
rect 12572 61794 12628 63868
rect 12684 62468 12740 65996
rect 12796 65958 12852 65996
rect 12908 67060 12964 67070
rect 12908 65828 12964 67004
rect 12796 65772 12964 65828
rect 13020 66050 13076 66062
rect 13020 65998 13022 66050
rect 13074 65998 13076 66050
rect 12796 62916 12852 65772
rect 13020 65492 13076 65998
rect 13020 65426 13076 65436
rect 12908 64708 12964 64718
rect 13132 64708 13188 74620
rect 13356 74228 13412 74732
rect 13356 74162 13412 74172
rect 13356 73108 13412 73118
rect 13244 73106 13412 73108
rect 13244 73054 13358 73106
rect 13410 73054 13412 73106
rect 13244 73052 13412 73054
rect 13244 72324 13300 73052
rect 13356 73042 13412 73052
rect 13244 71204 13300 72268
rect 13468 71764 13524 75852
rect 13580 75682 13636 76300
rect 13804 76354 13860 77308
rect 13804 76302 13806 76354
rect 13858 76302 13860 76354
rect 13804 76020 13860 76302
rect 13804 75954 13860 75964
rect 13580 75630 13582 75682
rect 13634 75630 13636 75682
rect 13580 75618 13636 75630
rect 13916 75908 13972 75918
rect 13692 75572 13748 75582
rect 13692 75348 13748 75516
rect 13916 75570 13972 75852
rect 13916 75518 13918 75570
rect 13970 75518 13972 75570
rect 13916 75506 13972 75518
rect 14028 75684 14084 75694
rect 13804 75460 13860 75470
rect 13804 75366 13860 75404
rect 13692 73948 13748 75292
rect 14028 75012 14084 75628
rect 13916 74956 14084 75012
rect 13804 74116 13860 74126
rect 13916 74116 13972 74956
rect 14028 74788 14084 74798
rect 14028 74786 14308 74788
rect 14028 74734 14030 74786
rect 14082 74734 14308 74786
rect 14028 74732 14308 74734
rect 14028 74722 14084 74732
rect 13804 74114 13972 74116
rect 13804 74062 13806 74114
rect 13858 74062 13972 74114
rect 13804 74060 13972 74062
rect 13804 74050 13860 74060
rect 13468 71698 13524 71708
rect 13580 73892 13748 73948
rect 13916 73948 13972 74060
rect 14140 74116 14196 74126
rect 13916 73892 14084 73948
rect 13244 71138 13300 71148
rect 13356 71652 13412 71662
rect 13356 68292 13412 71596
rect 13468 71540 13524 71550
rect 13468 70588 13524 71484
rect 13580 71316 13636 73892
rect 14028 73330 14084 73892
rect 14028 73278 14030 73330
rect 14082 73278 14084 73330
rect 13692 72434 13748 72446
rect 13692 72382 13694 72434
rect 13746 72382 13748 72434
rect 13692 71540 13748 72382
rect 13692 71474 13748 71484
rect 13804 72322 13860 72334
rect 13804 72270 13806 72322
rect 13858 72270 13860 72322
rect 13804 71988 13860 72270
rect 13580 71250 13636 71260
rect 13804 71092 13860 71932
rect 14028 71652 14084 73278
rect 14028 71586 14084 71596
rect 13916 71316 13972 71326
rect 14140 71316 14196 74060
rect 14252 72772 14308 74732
rect 14252 72706 14308 72716
rect 14364 73892 14420 79884
rect 14476 79716 14532 79726
rect 14476 74226 14532 79660
rect 15148 79380 15204 79390
rect 14476 74174 14478 74226
rect 14530 74174 14532 74226
rect 14476 74162 14532 74174
rect 14588 77924 14644 77934
rect 14588 75794 14644 77868
rect 14588 75742 14590 75794
rect 14642 75742 14644 75794
rect 13916 71202 13972 71260
rect 13916 71150 13918 71202
rect 13970 71150 13972 71202
rect 13916 71138 13972 71150
rect 14028 71260 14196 71316
rect 14028 71204 14084 71260
rect 14364 71204 14420 73836
rect 14476 72322 14532 72334
rect 14476 72270 14478 72322
rect 14530 72270 14532 72322
rect 14476 71876 14532 72270
rect 14476 71810 14532 71820
rect 14364 71148 14532 71204
rect 13804 71026 13860 71036
rect 14028 70980 14084 71148
rect 14140 70980 14196 70990
rect 14364 70980 14420 70990
rect 14028 70978 14196 70980
rect 14028 70926 14142 70978
rect 14194 70926 14196 70978
rect 14028 70924 14196 70926
rect 14140 70914 14196 70924
rect 14252 70978 14420 70980
rect 14252 70926 14366 70978
rect 14418 70926 14420 70978
rect 14252 70924 14420 70926
rect 13692 70866 13748 70878
rect 13692 70814 13694 70866
rect 13746 70814 13748 70866
rect 13692 70756 13748 70814
rect 14252 70756 14308 70924
rect 14364 70914 14420 70924
rect 13468 70532 13636 70588
rect 13468 70194 13524 70206
rect 13468 70142 13470 70194
rect 13522 70142 13524 70194
rect 13468 69748 13524 70142
rect 13468 68964 13524 69692
rect 13468 68898 13524 68908
rect 12908 64036 12964 64652
rect 12908 63250 12964 63980
rect 12908 63198 12910 63250
rect 12962 63198 12964 63250
rect 12908 63186 12964 63198
rect 13020 64652 13188 64708
rect 13244 68236 13412 68292
rect 12796 62850 12852 62860
rect 13020 62692 13076 64652
rect 13020 62626 13076 62636
rect 13132 64148 13188 64158
rect 12684 62412 13076 62468
rect 12572 61742 12574 61794
rect 12626 61742 12628 61794
rect 12572 61730 12628 61742
rect 12684 62242 12740 62254
rect 12684 62190 12686 62242
rect 12738 62190 12740 62242
rect 12684 62130 12740 62190
rect 12684 62078 12686 62130
rect 12738 62078 12740 62130
rect 12684 61796 12740 62078
rect 12684 61730 12740 61740
rect 12908 62020 12964 62030
rect 12908 61794 12964 61964
rect 12908 61742 12910 61794
rect 12962 61742 12964 61794
rect 12908 61730 12964 61742
rect 12572 61572 12628 61582
rect 12460 61570 12628 61572
rect 12460 61518 12574 61570
rect 12626 61518 12628 61570
rect 12460 61516 12628 61518
rect 12348 60674 12404 61516
rect 12572 61506 12628 61516
rect 13020 60900 13076 62412
rect 12348 60622 12350 60674
rect 12402 60622 12404 60674
rect 12348 60564 12404 60622
rect 12348 60498 12404 60508
rect 12460 60844 13076 60900
rect 12124 60274 12180 60284
rect 12012 59780 12068 60172
rect 11676 59724 12068 59780
rect 11676 59442 11732 59724
rect 11676 59390 11678 59442
rect 11730 59390 11732 59442
rect 11676 59378 11732 59390
rect 12460 59442 12516 60844
rect 12796 60674 12852 60686
rect 12796 60622 12798 60674
rect 12850 60622 12852 60674
rect 12684 60564 12740 60574
rect 12684 60114 12740 60508
rect 12684 60062 12686 60114
rect 12738 60062 12740 60114
rect 12684 60050 12740 60062
rect 12796 60116 12852 60622
rect 12796 59668 12852 60060
rect 13020 60564 13076 60574
rect 12796 59602 12852 59612
rect 12908 59780 12964 59790
rect 12460 59390 12462 59442
rect 12514 59390 12516 59442
rect 12460 59378 12516 59390
rect 11676 58548 11732 58558
rect 11564 58546 11732 58548
rect 11564 58494 11678 58546
rect 11730 58494 11732 58546
rect 11564 58492 11732 58494
rect 11228 58482 11284 58492
rect 11676 58482 11732 58492
rect 12124 58548 12180 58558
rect 12124 58454 12180 58492
rect 12572 58548 12628 58558
rect 12572 58454 12628 58492
rect 12012 58212 12068 58222
rect 11564 57876 11620 57886
rect 11116 57874 11564 57876
rect 11116 57822 11118 57874
rect 11170 57822 11564 57874
rect 11116 57820 11564 57822
rect 10444 57810 10500 57820
rect 11116 57810 11172 57820
rect 11564 57744 11620 57820
rect 12012 57874 12068 58156
rect 12012 57822 12014 57874
rect 12066 57822 12068 57874
rect 12012 57810 12068 57822
rect 12460 57876 12516 57886
rect 12908 57876 12964 59724
rect 13020 59442 13076 60508
rect 13020 59390 13022 59442
rect 13074 59390 13076 59442
rect 13020 59378 13076 59390
rect 13020 58548 13076 58558
rect 13132 58548 13188 64092
rect 13020 58546 13188 58548
rect 13020 58494 13022 58546
rect 13074 58494 13188 58546
rect 13020 58492 13188 58494
rect 13020 58482 13076 58492
rect 13020 57876 13076 57886
rect 12908 57874 13076 57876
rect 12908 57822 13022 57874
rect 13074 57822 13076 57874
rect 12908 57820 13076 57822
rect 12460 57782 12516 57820
rect 13020 57810 13076 57820
rect 12460 57652 12516 57662
rect 10332 51986 10388 51996
rect 11676 56644 11732 56654
rect 11676 50372 11732 56588
rect 11676 50306 11732 50316
rect 8204 5842 8260 5852
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 7308 4450 7364 4462
rect 7308 4398 7310 4450
rect 7362 4398 7364 4450
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6972 3668 7028 3678
rect 3500 3556 3556 3566
rect 3500 3462 3556 3500
rect 4284 3556 4340 3566
rect 4284 3462 4340 3500
rect 2604 3444 2660 3454
rect 2268 3442 2660 3444
rect 2268 3390 2606 3442
rect 2658 3390 2660 3442
rect 2268 3388 2660 3390
rect 2268 800 2324 3388
rect 2604 3378 2660 3388
rect 6972 800 7028 3612
rect 7308 3554 7364 4398
rect 9996 4452 10052 48300
rect 11004 6132 11060 6142
rect 11004 5906 11060 6076
rect 12460 6132 12516 57596
rect 13244 57540 13300 68236
rect 13468 65378 13524 65390
rect 13468 65326 13470 65378
rect 13522 65326 13524 65378
rect 13468 64820 13524 65326
rect 13580 64932 13636 70532
rect 13692 70308 13748 70700
rect 14028 70700 14308 70756
rect 14028 70588 14084 70700
rect 14476 70588 14532 71148
rect 14588 70756 14644 75742
rect 15148 74452 15204 79324
rect 15904 79200 16016 80000
rect 17948 79492 18004 79502
rect 15932 78820 15988 79200
rect 15932 77700 15988 78764
rect 17388 78932 17444 78942
rect 15932 77644 16100 77700
rect 15932 76354 15988 76366
rect 15932 76302 15934 76354
rect 15986 76302 15988 76354
rect 15932 76244 15988 76302
rect 15932 76178 15988 76188
rect 14812 73556 14868 73566
rect 14812 73442 14868 73500
rect 14812 73390 14814 73442
rect 14866 73390 14868 73442
rect 14812 73378 14868 73390
rect 15036 72436 15092 72446
rect 14588 70690 14644 70700
rect 14812 70754 14868 70766
rect 14812 70702 14814 70754
rect 14866 70702 14868 70754
rect 13692 70242 13748 70252
rect 13916 70532 14084 70588
rect 14364 70532 14532 70588
rect 13692 69522 13748 69534
rect 13692 69470 13694 69522
rect 13746 69470 13748 69522
rect 13692 69412 13748 69470
rect 13692 69346 13748 69356
rect 13804 67954 13860 67966
rect 13804 67902 13806 67954
rect 13858 67902 13860 67954
rect 13804 67844 13860 67902
rect 13804 67778 13860 67788
rect 13692 66388 13748 66398
rect 13692 66294 13748 66332
rect 13804 65490 13860 65502
rect 13804 65438 13806 65490
rect 13858 65438 13860 65490
rect 13804 65380 13860 65438
rect 13804 65314 13860 65324
rect 13580 64866 13636 64876
rect 13468 64754 13524 64764
rect 13916 64708 13972 70532
rect 14252 70084 14308 70094
rect 14140 70082 14308 70084
rect 14140 70030 14254 70082
rect 14306 70030 14308 70082
rect 14140 70028 14308 70030
rect 13916 64484 13972 64652
rect 13580 64260 13636 64270
rect 13580 63922 13636 64204
rect 13580 63870 13582 63922
rect 13634 63870 13636 63922
rect 13356 62804 13412 62814
rect 13356 62578 13412 62748
rect 13356 62526 13358 62578
rect 13410 62526 13412 62578
rect 13356 62468 13412 62526
rect 13356 62402 13412 62412
rect 13468 62580 13524 62590
rect 13580 62580 13636 63870
rect 13692 64148 13748 64158
rect 13692 63698 13748 64092
rect 13916 63810 13972 64428
rect 14028 68068 14084 68078
rect 14028 64818 14084 68012
rect 14028 64766 14030 64818
rect 14082 64766 14084 64818
rect 14028 64148 14084 64766
rect 14028 64082 14084 64092
rect 13916 63758 13918 63810
rect 13970 63758 13972 63810
rect 13916 63746 13972 63758
rect 13692 63646 13694 63698
rect 13746 63646 13748 63698
rect 13692 63634 13748 63646
rect 14140 63588 14196 70028
rect 14252 70018 14308 70028
rect 14252 67842 14308 67854
rect 14252 67790 14254 67842
rect 14306 67790 14308 67842
rect 14252 67060 14308 67790
rect 14364 67618 14420 70532
rect 14812 68180 14868 70702
rect 14476 68124 14868 68180
rect 14924 70644 14980 70654
rect 14476 67842 14532 68124
rect 14476 67790 14478 67842
rect 14530 67790 14532 67842
rect 14476 67778 14532 67790
rect 14812 67844 14868 67854
rect 14364 67566 14366 67618
rect 14418 67566 14420 67618
rect 14364 67554 14420 67566
rect 14252 66994 14308 67004
rect 14476 67060 14532 67070
rect 14364 66948 14420 66958
rect 14364 66854 14420 66892
rect 14476 66612 14532 67004
rect 14588 66612 14644 66622
rect 14476 66556 14588 66612
rect 14588 66546 14644 66556
rect 14364 66164 14420 66174
rect 14252 64932 14308 64942
rect 14252 64838 14308 64876
rect 14364 64706 14420 66108
rect 14812 66164 14868 67788
rect 14924 67170 14980 70588
rect 14924 67118 14926 67170
rect 14978 67118 14980 67170
rect 14924 67106 14980 67118
rect 15036 66388 15092 72380
rect 15148 68852 15204 74396
rect 15484 76020 15540 76030
rect 15372 71204 15428 71214
rect 15260 70978 15316 70990
rect 15260 70926 15262 70978
rect 15314 70926 15316 70978
rect 15260 70868 15316 70926
rect 15260 70802 15316 70812
rect 15148 68786 15204 68796
rect 15372 70644 15428 71148
rect 15372 67172 15428 70588
rect 15260 67116 15428 67172
rect 15148 67060 15204 67070
rect 15148 66966 15204 67004
rect 15260 66836 15316 67116
rect 15372 66948 15428 66958
rect 15484 66948 15540 75964
rect 16044 75012 16100 77644
rect 16716 76468 16772 76478
rect 16716 76374 16772 76412
rect 16828 75796 16884 75806
rect 16828 75702 16884 75740
rect 16044 74946 16100 74956
rect 16940 75684 16996 75694
rect 16940 74900 16996 75628
rect 17388 75012 17444 78876
rect 17724 76466 17780 76478
rect 17724 76414 17726 76466
rect 17778 76414 17780 76466
rect 17500 75684 17556 75694
rect 17724 75684 17780 76414
rect 17556 75628 17780 75684
rect 17500 75590 17556 75628
rect 17724 75124 17780 75134
rect 17388 74956 17556 75012
rect 16940 74898 17444 74900
rect 16940 74846 16942 74898
rect 16994 74846 17444 74898
rect 16940 74844 17444 74846
rect 16940 74834 16996 74844
rect 16156 74786 16212 74798
rect 16156 74734 16158 74786
rect 16210 74734 16212 74786
rect 16156 69972 16212 74734
rect 16604 74340 16660 74350
rect 16604 74226 16660 74284
rect 16604 74174 16606 74226
rect 16658 74174 16660 74226
rect 16604 74162 16660 74174
rect 17164 74114 17220 74126
rect 17164 74062 17166 74114
rect 17218 74062 17220 74114
rect 16940 73218 16996 73230
rect 16940 73166 16942 73218
rect 16994 73166 16996 73218
rect 16716 72436 16772 72446
rect 16716 72342 16772 72380
rect 16716 71762 16772 71774
rect 16716 71710 16718 71762
rect 16770 71710 16772 71762
rect 16380 70644 16436 70654
rect 16380 70082 16436 70588
rect 16716 70644 16772 71710
rect 16380 70030 16382 70082
rect 16434 70030 16436 70082
rect 16380 70018 16436 70030
rect 16492 70532 16548 70542
rect 16156 69906 16212 69916
rect 15820 69298 15876 69310
rect 15820 69246 15822 69298
rect 15874 69246 15876 69298
rect 15596 68404 15652 68414
rect 15596 67842 15652 68348
rect 15708 67956 15764 67966
rect 15708 67862 15764 67900
rect 15596 67790 15598 67842
rect 15650 67790 15652 67842
rect 15596 67396 15652 67790
rect 15596 67330 15652 67340
rect 15708 67730 15764 67742
rect 15708 67678 15710 67730
rect 15762 67678 15764 67730
rect 15596 67060 15652 67070
rect 15596 66966 15652 67004
rect 15372 66946 15540 66948
rect 15372 66894 15374 66946
rect 15426 66894 15540 66946
rect 15372 66892 15540 66894
rect 15372 66882 15428 66892
rect 14812 66098 14868 66108
rect 14924 66332 15036 66388
rect 14812 65492 14868 65502
rect 14812 65398 14868 65436
rect 14364 64654 14366 64706
rect 14418 64654 14420 64706
rect 14364 64642 14420 64654
rect 14924 64148 14980 66332
rect 15036 66322 15092 66332
rect 15148 66780 15316 66836
rect 14028 63532 14196 63588
rect 14812 64092 14980 64148
rect 15036 64708 15092 64718
rect 15036 64146 15092 64652
rect 15148 64372 15204 66780
rect 15708 66276 15764 67678
rect 15820 67284 15876 69246
rect 16492 68964 16548 70476
rect 16604 69748 16660 69758
rect 16604 69410 16660 69692
rect 16604 69358 16606 69410
rect 16658 69358 16660 69410
rect 16604 69346 16660 69358
rect 16380 68292 16436 68302
rect 16268 67844 16324 67854
rect 16268 67750 16324 67788
rect 15820 67218 15876 67228
rect 15932 67620 15988 67630
rect 15708 66210 15764 66220
rect 15820 66162 15876 66174
rect 15820 66110 15822 66162
rect 15874 66110 15876 66162
rect 15820 65828 15876 66110
rect 15820 65762 15876 65772
rect 15596 65492 15652 65502
rect 15596 65398 15652 65436
rect 15932 65044 15988 67564
rect 16044 66836 16100 66846
rect 16044 66834 16212 66836
rect 16044 66782 16046 66834
rect 16098 66782 16212 66834
rect 16044 66780 16212 66782
rect 16044 66770 16100 66780
rect 15932 64978 15988 64988
rect 16044 66052 16100 66062
rect 15372 64932 15428 64942
rect 15372 64838 15428 64876
rect 16044 64930 16100 65996
rect 16044 64878 16046 64930
rect 16098 64878 16100 64930
rect 15484 64708 15540 64718
rect 15484 64706 15652 64708
rect 15484 64654 15486 64706
rect 15538 64654 15652 64706
rect 15484 64652 15652 64654
rect 15484 64642 15540 64652
rect 15148 64316 15316 64372
rect 15260 64260 15316 64316
rect 15036 64094 15038 64146
rect 15090 64094 15092 64146
rect 13804 63138 13860 63150
rect 13804 63086 13806 63138
rect 13858 63086 13860 63138
rect 13692 63028 13748 63038
rect 13692 62934 13748 62972
rect 13468 62578 13636 62580
rect 13468 62526 13470 62578
rect 13522 62526 13636 62578
rect 13468 62524 13636 62526
rect 13692 62804 13748 62814
rect 13692 62578 13748 62748
rect 13692 62526 13694 62578
rect 13746 62526 13748 62578
rect 13356 61796 13412 61806
rect 13356 60898 13412 61740
rect 13356 60846 13358 60898
rect 13410 60846 13412 60898
rect 13356 60116 13412 60846
rect 13468 61010 13524 62524
rect 13692 62514 13748 62526
rect 13580 62356 13636 62366
rect 13580 62262 13636 62300
rect 13804 62188 13860 63086
rect 13692 62132 13860 62188
rect 13916 62354 13972 62366
rect 13916 62302 13918 62354
rect 13970 62302 13972 62354
rect 13692 62020 13748 62132
rect 13692 61954 13748 61964
rect 13804 61908 13860 61918
rect 13804 61682 13860 61852
rect 13804 61630 13806 61682
rect 13858 61630 13860 61682
rect 13804 61618 13860 61630
rect 13916 61684 13972 62302
rect 14028 62244 14084 63532
rect 14364 63140 14420 63150
rect 14364 63046 14420 63084
rect 14028 62178 14084 62188
rect 14364 62242 14420 62254
rect 14364 62190 14366 62242
rect 14418 62190 14420 62242
rect 14364 62132 14420 62190
rect 14252 62076 14364 62132
rect 13916 61618 13972 61628
rect 14140 61908 14196 61918
rect 13692 61348 13748 61358
rect 13692 61254 13748 61292
rect 13916 61346 13972 61358
rect 13916 61294 13918 61346
rect 13970 61294 13972 61346
rect 13916 61236 13972 61294
rect 13468 60958 13470 61010
rect 13522 60958 13524 61010
rect 13468 60900 13524 60958
rect 13692 61012 13748 61022
rect 13692 60918 13748 60956
rect 13468 60834 13524 60844
rect 13916 60564 13972 61180
rect 14028 60900 14084 60910
rect 14028 60806 14084 60844
rect 13916 60498 13972 60508
rect 14140 60228 14196 61852
rect 14252 61124 14308 62076
rect 14364 62066 14420 62076
rect 14364 61908 14420 61918
rect 14364 61570 14420 61852
rect 14364 61518 14366 61570
rect 14418 61518 14420 61570
rect 14364 61506 14420 61518
rect 14700 61460 14756 61470
rect 14700 61366 14756 61404
rect 14252 61058 14308 61068
rect 14364 61348 14420 61358
rect 14364 61012 14420 61292
rect 14476 61012 14532 61022
rect 14364 61010 14532 61012
rect 14364 60958 14478 61010
rect 14530 60958 14532 61010
rect 14364 60956 14532 60958
rect 14476 60946 14532 60956
rect 13580 60116 13636 60126
rect 13412 60114 13636 60116
rect 13412 60062 13582 60114
rect 13634 60062 13636 60114
rect 13412 60060 13636 60062
rect 13356 59984 13412 60060
rect 13580 60050 13636 60060
rect 13580 59332 13636 59342
rect 13580 59238 13636 59276
rect 14028 59106 14084 59118
rect 14028 59054 14030 59106
rect 14082 59054 14084 59106
rect 13692 58548 13748 58558
rect 13692 58454 13748 58492
rect 14028 58210 14084 59054
rect 14028 58158 14030 58210
rect 14082 58158 14084 58210
rect 13804 57764 13860 57774
rect 13356 57540 13412 57550
rect 13244 57484 13356 57540
rect 13356 57446 13412 57484
rect 13580 56868 13636 56878
rect 13580 56774 13636 56812
rect 12572 56642 12628 56654
rect 12572 56590 12574 56642
rect 12626 56590 12628 56642
rect 12572 56532 12628 56590
rect 12908 56644 12964 56654
rect 12908 56550 12964 56588
rect 12572 56466 12628 56476
rect 13804 36708 13860 57708
rect 14028 57540 14084 58158
rect 14028 57474 14084 57484
rect 14140 56978 14196 60172
rect 14252 60900 14308 60910
rect 14252 60116 14308 60844
rect 14700 60116 14756 60126
rect 14252 60114 14756 60116
rect 14252 60062 14254 60114
rect 14306 60062 14702 60114
rect 14754 60062 14756 60114
rect 14252 60060 14756 60062
rect 14252 60050 14308 60060
rect 14700 60050 14756 60060
rect 14812 58548 14868 64092
rect 15036 62578 15092 64094
rect 15148 64148 15204 64158
rect 15148 64054 15204 64092
rect 15260 64146 15316 64204
rect 15260 64094 15262 64146
rect 15314 64094 15316 64146
rect 15260 63476 15316 64094
rect 15484 63924 15540 63934
rect 15484 63830 15540 63868
rect 15260 63410 15316 63420
rect 15260 63252 15316 63262
rect 15260 63028 15316 63196
rect 15596 63140 15652 64652
rect 15708 64706 15764 64718
rect 15708 64654 15710 64706
rect 15762 64654 15764 64706
rect 15708 64036 15764 64654
rect 15708 63970 15764 63980
rect 15932 64708 15988 64718
rect 15708 63698 15764 63710
rect 15708 63646 15710 63698
rect 15762 63646 15764 63698
rect 15708 63252 15764 63646
rect 15932 63362 15988 64652
rect 16044 64484 16100 64878
rect 16044 64418 16100 64428
rect 15932 63310 15934 63362
rect 15986 63310 15988 63362
rect 15932 63298 15988 63310
rect 16044 63476 16100 63486
rect 15708 63186 15764 63196
rect 16044 63250 16100 63420
rect 16044 63198 16046 63250
rect 16098 63198 16100 63250
rect 15596 63074 15652 63084
rect 15260 62962 15316 62972
rect 15596 62692 15652 62702
rect 15036 62526 15038 62578
rect 15090 62526 15092 62578
rect 14924 62354 14980 62366
rect 14924 62302 14926 62354
rect 14978 62302 14980 62354
rect 14924 61460 14980 62302
rect 15036 62188 15092 62526
rect 15260 62580 15316 62590
rect 15260 62486 15316 62524
rect 15036 62132 15316 62188
rect 14924 61394 14980 61404
rect 15036 61684 15092 61694
rect 15036 61010 15092 61628
rect 15148 61572 15204 61582
rect 15148 61478 15204 61516
rect 15036 60958 15038 61010
rect 15090 60958 15092 61010
rect 14924 60900 14980 60910
rect 14924 59442 14980 60844
rect 15036 60788 15092 60958
rect 15260 61012 15316 62132
rect 15372 61012 15428 61022
rect 15260 61010 15428 61012
rect 15260 60958 15374 61010
rect 15426 60958 15428 61010
rect 15260 60956 15428 60958
rect 15372 60946 15428 60956
rect 15036 60722 15092 60732
rect 15372 59892 15428 59902
rect 15372 59798 15428 59836
rect 14924 59390 14926 59442
rect 14978 59390 14980 59442
rect 14924 59378 14980 59390
rect 15484 59444 15540 59454
rect 15484 59350 15540 59388
rect 15596 58658 15652 62636
rect 15820 62692 15876 62702
rect 15820 62578 15876 62636
rect 15820 62526 15822 62578
rect 15874 62526 15876 62578
rect 15820 62514 15876 62526
rect 15932 62466 15988 62478
rect 15932 62414 15934 62466
rect 15986 62414 15988 62466
rect 15708 62132 15764 62142
rect 15708 62038 15764 62076
rect 15932 62020 15988 62414
rect 16044 62132 16100 63198
rect 16044 62066 16100 62076
rect 15932 61954 15988 61964
rect 15596 58606 15598 58658
rect 15650 58606 15652 58658
rect 15596 58594 15652 58606
rect 15708 61796 15764 61806
rect 15036 58548 15092 58558
rect 15372 58548 15428 58558
rect 14812 58546 15092 58548
rect 14812 58494 15038 58546
rect 15090 58494 15092 58546
rect 14812 58492 15092 58494
rect 15036 58482 15092 58492
rect 15148 58492 15372 58548
rect 14476 58212 14532 58222
rect 14252 57652 14308 57662
rect 14252 57558 14308 57596
rect 14140 56926 14142 56978
rect 14194 56926 14196 56978
rect 14140 56914 14196 56926
rect 14476 56308 14532 58156
rect 14700 57876 14756 57886
rect 14700 57540 14756 57820
rect 15148 57876 15204 58492
rect 15372 58454 15428 58492
rect 15148 57744 15204 57820
rect 14700 57446 14756 57484
rect 14476 56242 14532 56252
rect 15148 56868 15204 56878
rect 15148 41860 15204 56812
rect 15708 55076 15764 61740
rect 16156 61794 16212 66780
rect 16380 65714 16436 68236
rect 16492 66274 16548 68908
rect 16604 69188 16660 69198
rect 16604 67730 16660 69132
rect 16716 68626 16772 70588
rect 16716 68574 16718 68626
rect 16770 68574 16772 68626
rect 16716 68562 16772 68574
rect 16940 70532 16996 73166
rect 16604 67678 16606 67730
rect 16658 67678 16660 67730
rect 16604 67666 16660 67678
rect 16716 67732 16772 67742
rect 16604 67060 16660 67098
rect 16604 66994 16660 67004
rect 16604 66834 16660 66846
rect 16604 66782 16606 66834
rect 16658 66782 16660 66834
rect 16604 66724 16660 66782
rect 16604 66658 16660 66668
rect 16492 66222 16494 66274
rect 16546 66222 16548 66274
rect 16492 66210 16548 66222
rect 16716 65828 16772 67676
rect 16828 67284 16884 67294
rect 16828 65940 16884 67228
rect 16940 67172 16996 70476
rect 17164 69748 17220 74062
rect 17388 72546 17444 74844
rect 17388 72494 17390 72546
rect 17442 72494 17444 72546
rect 17388 72482 17444 72494
rect 17500 74788 17556 74956
rect 17164 69682 17220 69692
rect 17388 71876 17444 71886
rect 17388 70084 17444 71820
rect 17164 69524 17220 69534
rect 16940 67106 16996 67116
rect 17052 69522 17220 69524
rect 17052 69470 17166 69522
rect 17218 69470 17220 69522
rect 17052 69468 17220 69470
rect 16940 66948 16996 66958
rect 16940 66854 16996 66892
rect 16828 65884 16996 65940
rect 16380 65662 16382 65714
rect 16434 65662 16436 65714
rect 16380 65650 16436 65662
rect 16492 65772 16772 65828
rect 16268 65604 16324 65614
rect 16268 65510 16324 65548
rect 16492 65492 16548 65772
rect 16380 65436 16548 65492
rect 16604 65492 16660 65502
rect 16268 65380 16324 65390
rect 16268 65286 16324 65324
rect 16380 64596 16436 65436
rect 16604 65398 16660 65436
rect 16716 65490 16772 65502
rect 16716 65438 16718 65490
rect 16770 65438 16772 65490
rect 16716 65268 16772 65438
rect 16716 65202 16772 65212
rect 16380 64146 16436 64540
rect 16380 64094 16382 64146
rect 16434 64094 16436 64146
rect 16380 64082 16436 64094
rect 16492 65044 16548 65054
rect 16492 64146 16548 64988
rect 16828 64706 16884 64718
rect 16828 64654 16830 64706
rect 16882 64654 16884 64706
rect 16492 64094 16494 64146
rect 16546 64094 16548 64146
rect 16492 64082 16548 64094
rect 16604 64484 16660 64494
rect 16604 64148 16660 64428
rect 16828 64148 16884 64654
rect 16940 64260 16996 65884
rect 17052 65828 17108 69468
rect 17164 69458 17220 69468
rect 17164 67956 17220 67966
rect 17164 67862 17220 67900
rect 17388 66948 17444 70028
rect 17500 67284 17556 74732
rect 17724 74788 17780 75068
rect 17724 74786 17892 74788
rect 17724 74734 17726 74786
rect 17778 74734 17892 74786
rect 17724 74732 17892 74734
rect 17724 74722 17780 74732
rect 17724 73332 17780 73342
rect 17836 73332 17892 74732
rect 17948 74226 18004 79436
rect 20272 79200 20384 80000
rect 24640 79200 24752 80000
rect 28812 79716 28868 79726
rect 28364 79604 28420 79614
rect 28420 79548 28644 79604
rect 28364 79538 28420 79548
rect 18396 79156 18452 79166
rect 17948 74174 17950 74226
rect 18002 74174 18004 74226
rect 17948 74162 18004 74174
rect 18060 76132 18116 76142
rect 17948 73332 18004 73342
rect 17836 73330 18004 73332
rect 17836 73278 17950 73330
rect 18002 73278 18004 73330
rect 17836 73276 18004 73278
rect 18060 73332 18116 76076
rect 18396 75684 18452 79100
rect 18732 79044 18788 79054
rect 18508 76356 18564 76366
rect 18508 76262 18564 76300
rect 18620 75908 18676 75918
rect 18396 75628 18564 75684
rect 18172 75458 18228 75470
rect 18172 75406 18174 75458
rect 18226 75406 18228 75458
rect 18172 75348 18228 75406
rect 18172 75282 18228 75292
rect 18284 75458 18340 75470
rect 18284 75406 18286 75458
rect 18338 75406 18340 75458
rect 18172 73332 18228 73342
rect 18060 73330 18228 73332
rect 18060 73278 18174 73330
rect 18226 73278 18228 73330
rect 18060 73276 18228 73278
rect 17724 73238 17780 73276
rect 17948 73266 18004 73276
rect 17724 73108 17780 73118
rect 17612 70756 17668 70766
rect 17612 70082 17668 70700
rect 17612 70030 17614 70082
rect 17666 70030 17668 70082
rect 17612 70018 17668 70030
rect 17724 67620 17780 73052
rect 18172 72660 18228 73276
rect 18284 72772 18340 75406
rect 18396 75460 18452 75470
rect 18396 74564 18452 75404
rect 18396 74498 18452 74508
rect 18508 74340 18564 75628
rect 18620 75570 18676 75852
rect 18620 75518 18622 75570
rect 18674 75518 18676 75570
rect 18620 75506 18676 75518
rect 18732 75236 18788 78988
rect 20300 78596 20356 79200
rect 20412 78596 20468 78606
rect 20300 78540 20412 78596
rect 20188 78148 20244 78158
rect 19068 78036 19124 78046
rect 18620 75180 18788 75236
rect 18844 76580 18900 76590
rect 18620 74788 18676 75180
rect 18732 75012 18788 75022
rect 18732 74918 18788 74956
rect 18620 74732 18788 74788
rect 18396 74284 18564 74340
rect 18620 74564 18676 74574
rect 18396 73108 18452 74284
rect 18508 73444 18564 73454
rect 18508 73350 18564 73388
rect 18396 73014 18452 73052
rect 18284 72716 18452 72772
rect 18172 72604 18340 72660
rect 18284 72546 18340 72604
rect 18284 72494 18286 72546
rect 18338 72494 18340 72546
rect 18284 72482 18340 72494
rect 18396 72548 18452 72716
rect 18396 72482 18452 72492
rect 18508 72548 18564 72558
rect 18620 72548 18676 74508
rect 18508 72546 18676 72548
rect 18508 72494 18510 72546
rect 18562 72494 18676 72546
rect 18508 72492 18676 72494
rect 18508 72482 18564 72492
rect 18060 72436 18116 72446
rect 17948 72434 18116 72436
rect 17948 72382 18062 72434
rect 18114 72382 18116 72434
rect 17948 72380 18116 72382
rect 17948 70588 18004 72380
rect 18060 72370 18116 72380
rect 18172 72436 18228 72446
rect 18060 71988 18116 71998
rect 18172 71988 18228 72380
rect 18396 72322 18452 72334
rect 18396 72270 18398 72322
rect 18450 72270 18452 72322
rect 18284 71988 18340 71998
rect 18172 71986 18340 71988
rect 18172 71934 18286 71986
rect 18338 71934 18340 71986
rect 18172 71932 18340 71934
rect 18060 71894 18116 71932
rect 18284 71922 18340 71932
rect 18172 71652 18228 71662
rect 17836 70532 18004 70588
rect 18060 71650 18228 71652
rect 18060 71598 18174 71650
rect 18226 71598 18228 71650
rect 18060 71596 18228 71598
rect 17836 68740 17892 70532
rect 17948 70082 18004 70094
rect 17948 70030 17950 70082
rect 18002 70030 18004 70082
rect 17948 69860 18004 70030
rect 17948 69794 18004 69804
rect 18060 69076 18116 71596
rect 18172 71586 18228 71596
rect 18396 70980 18452 72270
rect 18396 70914 18452 70924
rect 18508 72324 18564 72334
rect 18172 70420 18228 70430
rect 18172 70418 18452 70420
rect 18172 70366 18174 70418
rect 18226 70366 18452 70418
rect 18172 70364 18452 70366
rect 18172 70354 18228 70364
rect 18172 70194 18228 70206
rect 18172 70142 18174 70194
rect 18226 70142 18228 70194
rect 18172 69636 18228 70142
rect 18396 70196 18452 70364
rect 18396 70130 18452 70140
rect 18508 70194 18564 72268
rect 18508 70142 18510 70194
rect 18562 70142 18564 70194
rect 18396 69972 18452 69982
rect 18172 69570 18228 69580
rect 18284 69860 18340 69870
rect 18060 69010 18116 69020
rect 17836 68674 17892 68684
rect 18172 68740 18228 68750
rect 18172 68626 18228 68684
rect 18172 68574 18174 68626
rect 18226 68574 18228 68626
rect 18172 68562 18228 68574
rect 18284 68628 18340 69804
rect 18396 68852 18452 69916
rect 18508 69636 18564 70142
rect 18508 69570 18564 69580
rect 18620 72324 18676 72334
rect 18732 72324 18788 74732
rect 18620 72322 18788 72324
rect 18620 72270 18622 72322
rect 18674 72270 18788 72322
rect 18620 72268 18788 72270
rect 18620 69412 18676 72268
rect 18732 71764 18788 71774
rect 18844 71764 18900 76524
rect 19068 73948 19124 77980
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19404 75794 19460 75806
rect 19404 75742 19406 75794
rect 19458 75742 19460 75794
rect 19404 75572 19460 75742
rect 19404 75506 19460 75516
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 20188 75012 20244 78092
rect 20132 74956 20244 75012
rect 20300 76468 20356 76478
rect 20300 75684 20356 76412
rect 19852 74788 19908 74798
rect 19628 74786 19908 74788
rect 19628 74734 19854 74786
rect 19906 74734 19908 74786
rect 19628 74732 19908 74734
rect 19068 73892 19348 73948
rect 19180 73444 19236 73454
rect 19068 73442 19236 73444
rect 19068 73390 19182 73442
rect 19234 73390 19236 73442
rect 19068 73388 19236 73390
rect 18732 71762 18900 71764
rect 18732 71710 18734 71762
rect 18786 71710 18900 71762
rect 18732 71708 18900 71710
rect 18956 72996 19012 73006
rect 18732 71652 18788 71708
rect 18732 71586 18788 71596
rect 18844 70532 18900 70542
rect 18844 70418 18900 70476
rect 18844 70366 18846 70418
rect 18898 70366 18900 70418
rect 18844 70354 18900 70366
rect 18620 69346 18676 69356
rect 18732 70194 18788 70206
rect 18732 70142 18734 70194
rect 18786 70142 18788 70194
rect 18508 68852 18564 68862
rect 18396 68850 18564 68852
rect 18396 68798 18510 68850
rect 18562 68798 18564 68850
rect 18396 68796 18564 68798
rect 18508 68786 18564 68796
rect 18396 68628 18452 68638
rect 18284 68626 18452 68628
rect 18284 68574 18398 68626
rect 18450 68574 18452 68626
rect 18284 68572 18452 68574
rect 18396 68562 18452 68572
rect 18508 68402 18564 68414
rect 18508 68350 18510 68402
rect 18562 68350 18564 68402
rect 18508 68292 18564 68350
rect 18508 68226 18564 68236
rect 17836 68068 17892 68078
rect 17836 67954 17892 68012
rect 17836 67902 17838 67954
rect 17890 67902 17892 67954
rect 17836 67890 17892 67902
rect 17724 67284 17780 67564
rect 18620 67844 18676 67854
rect 17500 67218 17556 67228
rect 17612 67228 17780 67284
rect 17948 67284 18004 67294
rect 17388 66882 17444 66892
rect 17612 66836 17668 67228
rect 17948 67190 18004 67228
rect 18284 67060 18340 67098
rect 18284 66994 18340 67004
rect 18508 67060 18564 67070
rect 18620 67060 18676 67788
rect 18732 67284 18788 70142
rect 18732 67218 18788 67228
rect 18844 70084 18900 70094
rect 18508 67058 18676 67060
rect 18508 67006 18510 67058
rect 18562 67006 18676 67058
rect 18508 67004 18676 67006
rect 18508 66994 18564 67004
rect 17836 66948 17892 66986
rect 18844 66948 18900 70028
rect 17836 66882 17892 66892
rect 18732 66892 18900 66948
rect 17612 66780 17780 66836
rect 17164 66612 17220 66622
rect 17164 66274 17220 66556
rect 17164 66222 17166 66274
rect 17218 66222 17220 66274
rect 17164 66210 17220 66222
rect 17388 66162 17444 66174
rect 17388 66110 17390 66162
rect 17442 66110 17444 66162
rect 17052 65772 17332 65828
rect 17164 64708 17220 64718
rect 17164 64614 17220 64652
rect 17164 64484 17220 64494
rect 16940 64204 17108 64260
rect 16604 64146 16772 64148
rect 16604 64094 16606 64146
rect 16658 64094 16772 64146
rect 16604 64092 16772 64094
rect 16604 64082 16660 64092
rect 16604 63700 16660 63710
rect 16380 63252 16436 63262
rect 16380 62580 16436 63196
rect 16492 62580 16548 62590
rect 16380 62578 16548 62580
rect 16380 62526 16494 62578
rect 16546 62526 16548 62578
rect 16380 62524 16548 62526
rect 16492 62514 16548 62524
rect 16604 62356 16660 63644
rect 16716 63364 16772 64092
rect 16828 64082 16884 64092
rect 17052 64036 17108 64204
rect 17052 63970 17108 63980
rect 16716 63298 16772 63308
rect 16940 63922 16996 63934
rect 16940 63870 16942 63922
rect 16994 63870 16996 63922
rect 16716 63138 16772 63150
rect 16716 63086 16718 63138
rect 16770 63086 16772 63138
rect 16716 63028 16772 63086
rect 16716 62962 16772 62972
rect 16716 62580 16772 62590
rect 16716 62486 16772 62524
rect 16492 62300 16660 62356
rect 16828 62354 16884 62366
rect 16828 62302 16830 62354
rect 16882 62302 16884 62354
rect 16156 61742 16158 61794
rect 16210 61742 16212 61794
rect 16156 61730 16212 61742
rect 16380 62020 16436 62030
rect 15820 61572 15876 61582
rect 15820 61478 15876 61516
rect 16044 61570 16100 61582
rect 16044 61518 16046 61570
rect 16098 61518 16100 61570
rect 16044 61460 16100 61518
rect 16044 61394 16100 61404
rect 15820 60900 15876 60910
rect 15820 60806 15876 60844
rect 16268 60676 16324 60686
rect 16380 60676 16436 61964
rect 16268 60674 16436 60676
rect 16268 60622 16270 60674
rect 16322 60622 16436 60674
rect 16268 60620 16436 60622
rect 16268 60228 16324 60620
rect 15820 60116 15876 60126
rect 16268 60116 16324 60172
rect 15820 60022 15876 60060
rect 16156 60060 16324 60116
rect 16380 60340 16436 60350
rect 16380 60114 16436 60284
rect 16380 60062 16382 60114
rect 16434 60062 16436 60114
rect 15932 59668 15988 59678
rect 15932 59442 15988 59612
rect 15932 59390 15934 59442
rect 15986 59390 15988 59442
rect 15932 59378 15988 59390
rect 15932 58772 15988 58782
rect 15932 58546 15988 58716
rect 15932 58494 15934 58546
rect 15986 58494 15988 58546
rect 15932 58482 15988 58494
rect 15708 55010 15764 55020
rect 16156 54964 16212 60060
rect 16380 60050 16436 60062
rect 16492 59442 16548 62300
rect 16828 62020 16884 62302
rect 16716 61460 16772 61470
rect 16716 61366 16772 61404
rect 16828 61012 16884 61964
rect 16940 61684 16996 63870
rect 16940 61348 16996 61628
rect 16940 61282 16996 61292
rect 17052 63812 17108 63822
rect 16828 60946 16884 60956
rect 17052 61010 17108 63756
rect 17164 62468 17220 64428
rect 17164 62402 17220 62412
rect 17164 62132 17220 62142
rect 17164 61682 17220 62076
rect 17276 61794 17332 65772
rect 17388 63700 17444 66110
rect 17500 66162 17556 66174
rect 17500 66110 17502 66162
rect 17554 66110 17556 66162
rect 17500 64932 17556 66110
rect 17724 65602 17780 66780
rect 18060 66834 18116 66846
rect 18060 66782 18062 66834
rect 18114 66782 18116 66834
rect 18060 66612 18116 66782
rect 18060 66546 18116 66556
rect 18284 66836 18340 66846
rect 18732 66836 18788 66892
rect 18284 66276 18340 66780
rect 18620 66780 18788 66836
rect 18508 66276 18564 66286
rect 18284 66274 18564 66276
rect 18284 66222 18510 66274
rect 18562 66222 18564 66274
rect 18284 66220 18564 66222
rect 18508 66210 18564 66220
rect 18620 66276 18676 66780
rect 18844 66724 18900 66734
rect 17724 65550 17726 65602
rect 17778 65550 17780 65602
rect 17724 65538 17780 65550
rect 17836 66164 17892 66174
rect 17500 64866 17556 64876
rect 17724 64820 17780 64830
rect 17836 64820 17892 66108
rect 18620 66162 18676 66220
rect 18620 66110 18622 66162
rect 18674 66110 18676 66162
rect 17948 66052 18004 66062
rect 17948 65958 18004 65996
rect 18620 65828 18676 66110
rect 18508 65772 18676 65828
rect 18732 66668 18844 66724
rect 18732 66500 18788 66668
rect 18844 66658 18900 66668
rect 17724 64818 17892 64820
rect 17724 64766 17726 64818
rect 17778 64766 17892 64818
rect 17724 64764 17892 64766
rect 17948 65716 18004 65726
rect 17948 65490 18004 65660
rect 18172 65716 18228 65726
rect 18172 65622 18228 65660
rect 17948 65438 17950 65490
rect 18002 65438 18004 65490
rect 17724 64754 17780 64764
rect 17948 64708 18004 65438
rect 18284 65490 18340 65502
rect 18284 65438 18286 65490
rect 18338 65438 18340 65490
rect 18172 65268 18228 65278
rect 17836 64652 18004 64708
rect 18060 65266 18228 65268
rect 18060 65214 18174 65266
rect 18226 65214 18228 65266
rect 18060 65212 18228 65214
rect 17388 63634 17444 63644
rect 17612 64484 17668 64494
rect 17612 63250 17668 64428
rect 17724 63812 17780 63822
rect 17724 63718 17780 63756
rect 17612 63198 17614 63250
rect 17666 63198 17668 63250
rect 17612 63186 17668 63198
rect 17500 63138 17556 63150
rect 17500 63086 17502 63138
rect 17554 63086 17556 63138
rect 17500 62020 17556 63086
rect 17612 63026 17668 63038
rect 17612 62974 17614 63026
rect 17666 62974 17668 63026
rect 17612 62580 17668 62974
rect 17612 62514 17668 62524
rect 17500 61954 17556 61964
rect 17276 61742 17278 61794
rect 17330 61742 17332 61794
rect 17276 61730 17332 61742
rect 17500 61794 17556 61806
rect 17500 61742 17502 61794
rect 17554 61742 17556 61794
rect 17164 61630 17166 61682
rect 17218 61630 17220 61682
rect 17164 61618 17220 61630
rect 17052 60958 17054 61010
rect 17106 60958 17108 61010
rect 17052 60946 17108 60958
rect 17500 61348 17556 61742
rect 17612 61348 17668 61358
rect 17500 61346 17668 61348
rect 17500 61294 17614 61346
rect 17666 61294 17668 61346
rect 17500 61292 17668 61294
rect 16828 60676 16884 60686
rect 16828 60114 16884 60620
rect 16828 60062 16830 60114
rect 16882 60062 16884 60114
rect 16828 60050 16884 60062
rect 17276 59780 17332 59790
rect 17276 59686 17332 59724
rect 16492 59390 16494 59442
rect 16546 59390 16548 59442
rect 16492 59378 16548 59390
rect 16940 59444 16996 59454
rect 16940 59350 16996 59388
rect 16828 58996 16884 59006
rect 16268 58658 16324 58670
rect 16268 58606 16270 58658
rect 16322 58606 16324 58658
rect 16268 58546 16324 58606
rect 16268 58494 16270 58546
rect 16322 58494 16324 58546
rect 16268 58482 16324 58494
rect 16716 58660 16772 58670
rect 16156 54898 16212 54908
rect 15148 40404 15204 41804
rect 15148 40338 15204 40348
rect 15932 40404 15988 40414
rect 13804 36642 13860 36652
rect 14812 6804 14868 6814
rect 12460 6000 12516 6076
rect 14364 6132 14420 6142
rect 14812 6132 14868 6748
rect 14364 6130 14868 6132
rect 14364 6078 14366 6130
rect 14418 6078 14814 6130
rect 14866 6078 14868 6130
rect 14364 6076 14868 6078
rect 14364 6066 14420 6076
rect 14812 6066 14868 6076
rect 15036 6020 15092 6030
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5842 11060 5854
rect 12124 5794 12180 5806
rect 12124 5742 12126 5794
rect 12178 5742 12180 5794
rect 11228 5682 11284 5694
rect 11228 5630 11230 5682
rect 11282 5630 11284 5682
rect 11228 4564 11284 5630
rect 11564 5682 11620 5694
rect 11564 5630 11566 5682
rect 11618 5630 11620 5682
rect 11452 5124 11508 5134
rect 11564 5124 11620 5630
rect 11452 5122 11620 5124
rect 11452 5070 11454 5122
rect 11506 5070 11620 5122
rect 11452 5068 11620 5070
rect 11452 5058 11508 5068
rect 11676 4900 11732 4910
rect 11228 4498 11284 4508
rect 11564 4898 11732 4900
rect 11564 4846 11678 4898
rect 11730 4846 11732 4898
rect 11564 4844 11732 4846
rect 9996 4386 10052 4396
rect 7644 4340 7700 4350
rect 7644 4246 7700 4284
rect 11340 4340 11396 4350
rect 11340 4246 11396 4284
rect 7868 3668 7924 3678
rect 7868 3574 7924 3612
rect 7308 3502 7310 3554
rect 7362 3502 7364 3554
rect 7308 3490 7364 3502
rect 11564 3554 11620 4844
rect 11676 4834 11732 4844
rect 11676 4564 11732 4574
rect 12124 4564 12180 5742
rect 12348 4564 12404 4574
rect 12124 4508 12348 4564
rect 11676 4338 11732 4508
rect 12348 4470 12404 4508
rect 14588 4564 14644 4574
rect 14588 4470 14644 4508
rect 11676 4286 11678 4338
rect 11730 4286 11732 4338
rect 11676 4274 11732 4286
rect 11900 4452 11956 4462
rect 11900 4338 11956 4396
rect 12796 4452 12852 4462
rect 12796 4358 12852 4396
rect 11900 4286 11902 4338
rect 11954 4286 11956 4338
rect 11900 4274 11956 4286
rect 15036 4340 15092 5964
rect 15932 6020 15988 40348
rect 15932 5954 15988 5964
rect 15372 5796 15428 5806
rect 15372 4564 15428 5740
rect 16716 5348 16772 58604
rect 16828 55300 16884 58940
rect 17164 58660 17220 58670
rect 17164 58546 17220 58604
rect 17164 58494 17166 58546
rect 17218 58494 17220 58546
rect 17164 58482 17220 58494
rect 17500 58436 17556 61292
rect 17612 61282 17668 61292
rect 17612 60900 17668 60910
rect 17612 60806 17668 60844
rect 17612 60116 17668 60126
rect 17836 60116 17892 64652
rect 18060 64148 18116 65212
rect 18172 65202 18228 65212
rect 18284 64820 18340 65438
rect 18508 65268 18564 65772
rect 18620 65604 18676 65614
rect 18732 65604 18788 66444
rect 18620 65602 18788 65604
rect 18620 65550 18622 65602
rect 18674 65550 18788 65602
rect 18620 65548 18788 65550
rect 18844 66050 18900 66062
rect 18844 65998 18846 66050
rect 18898 65998 18900 66050
rect 18620 65538 18676 65548
rect 18508 65212 18676 65268
rect 18284 64754 18340 64764
rect 18508 64708 18564 64718
rect 18396 64596 18452 64606
rect 18396 64502 18452 64540
rect 18284 64482 18340 64494
rect 18284 64430 18286 64482
rect 18338 64430 18340 64482
rect 17948 64092 18116 64148
rect 18172 64372 18228 64382
rect 18172 64146 18228 64316
rect 18172 64094 18174 64146
rect 18226 64094 18228 64146
rect 17948 62692 18004 64092
rect 18172 64082 18228 64094
rect 18284 64148 18340 64430
rect 18284 64082 18340 64092
rect 18508 64482 18564 64652
rect 18508 64430 18510 64482
rect 18562 64430 18564 64482
rect 17948 62626 18004 62636
rect 18060 63922 18116 63934
rect 18060 63870 18062 63922
rect 18114 63870 18116 63922
rect 17948 62242 18004 62254
rect 17948 62190 17950 62242
rect 18002 62190 18004 62242
rect 17948 61794 18004 62190
rect 17948 61742 17950 61794
rect 18002 61742 18004 61794
rect 17948 61730 18004 61742
rect 18060 61572 18116 63870
rect 18172 63924 18228 63934
rect 18396 63924 18452 63934
rect 18228 63868 18340 63924
rect 18172 63858 18228 63868
rect 18284 63810 18340 63868
rect 18396 63830 18452 63868
rect 18284 63758 18286 63810
rect 18338 63758 18340 63810
rect 18284 63746 18340 63758
rect 18508 63364 18564 64430
rect 18620 63700 18676 65212
rect 18620 63634 18676 63644
rect 18732 64372 18788 64382
rect 18396 63308 18564 63364
rect 18620 63364 18676 63374
rect 18396 63250 18452 63308
rect 18396 63198 18398 63250
rect 18450 63198 18452 63250
rect 18396 63186 18452 63198
rect 18620 63138 18676 63308
rect 18620 63086 18622 63138
rect 18674 63086 18676 63138
rect 18620 63074 18676 63086
rect 18060 61506 18116 61516
rect 18172 62356 18228 62366
rect 18172 62130 18228 62300
rect 18732 62188 18788 64316
rect 18844 64036 18900 65998
rect 18956 64932 19012 72940
rect 19068 65492 19124 73388
rect 19180 73378 19236 73388
rect 19180 71762 19236 71774
rect 19180 71710 19182 71762
rect 19234 71710 19236 71762
rect 19180 70866 19236 71710
rect 19180 70814 19182 70866
rect 19234 70814 19236 70866
rect 19180 70644 19236 70814
rect 19180 68626 19236 70588
rect 19292 69522 19348 73892
rect 19404 73330 19460 73342
rect 19404 73278 19406 73330
rect 19458 73278 19460 73330
rect 19404 72212 19460 73278
rect 19628 72548 19684 74732
rect 19852 74722 19908 74732
rect 20132 74676 20188 74956
rect 20300 74898 20356 75628
rect 20412 75570 20468 78540
rect 24556 78484 24612 78494
rect 22988 78372 23044 78382
rect 20636 76580 20692 76590
rect 20636 76354 20692 76524
rect 22316 76468 22372 76478
rect 20636 76302 20638 76354
rect 20690 76302 20692 76354
rect 20636 76290 20692 76302
rect 21420 76356 21476 76366
rect 21420 76262 21476 76300
rect 20412 75518 20414 75570
rect 20466 75518 20468 75570
rect 20412 75506 20468 75518
rect 21756 75682 21812 75694
rect 21756 75630 21758 75682
rect 21810 75630 21812 75682
rect 20300 74846 20302 74898
rect 20354 74846 20356 74898
rect 20132 74620 20244 74676
rect 20076 74228 20132 74238
rect 20076 74134 20132 74172
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 20188 73556 20244 74620
rect 20076 73500 20244 73556
rect 20076 73108 20132 73500
rect 20188 73332 20244 73342
rect 20300 73332 20356 74846
rect 21084 74788 21140 74798
rect 20188 73330 20356 73332
rect 20188 73278 20190 73330
rect 20242 73278 20356 73330
rect 20188 73276 20356 73278
rect 20412 74786 21140 74788
rect 20412 74734 21086 74786
rect 21138 74734 21140 74786
rect 20412 74732 21140 74734
rect 20188 73266 20244 73276
rect 20076 73052 20244 73108
rect 19740 72996 19796 73006
rect 19740 72770 19796 72940
rect 20188 72884 20244 73052
rect 20300 72884 20356 72894
rect 20188 72828 20300 72884
rect 19740 72718 19742 72770
rect 19794 72718 19796 72770
rect 19740 72706 19796 72718
rect 19628 72492 19796 72548
rect 19516 72324 19572 72334
rect 19516 72230 19572 72268
rect 19628 72322 19684 72334
rect 19628 72270 19630 72322
rect 19682 72270 19684 72322
rect 19404 70980 19460 72156
rect 19404 70914 19460 70924
rect 19516 70084 19572 70094
rect 19516 69990 19572 70028
rect 19628 69860 19684 72270
rect 19740 72324 19796 72492
rect 20300 72546 20356 72828
rect 20412 72658 20468 74732
rect 21084 74722 21140 74732
rect 21756 74676 21812 75630
rect 22316 75684 22372 76412
rect 22988 75794 23044 78316
rect 23548 77364 23604 77374
rect 23548 76578 23604 77308
rect 23548 76526 23550 76578
rect 23602 76526 23604 76578
rect 23548 76514 23604 76526
rect 24332 76468 24388 76478
rect 24332 76374 24388 76412
rect 22988 75742 22990 75794
rect 23042 75742 23044 75794
rect 22988 75730 23044 75742
rect 22316 75552 22372 75628
rect 24220 74898 24276 74910
rect 24220 74846 24222 74898
rect 24274 74846 24276 74898
rect 21532 74116 21588 74126
rect 20860 74004 20916 74014
rect 20860 74002 21028 74004
rect 20860 73950 20862 74002
rect 20914 73950 21028 74002
rect 20860 73948 21028 73950
rect 20860 73938 20916 73948
rect 20412 72606 20414 72658
rect 20466 72606 20468 72658
rect 20412 72594 20468 72606
rect 20524 73890 20580 73902
rect 20524 73838 20526 73890
rect 20578 73838 20580 73890
rect 20300 72494 20302 72546
rect 20354 72494 20356 72546
rect 20300 72482 20356 72494
rect 20412 72324 20468 72334
rect 19740 72268 20244 72324
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 20188 71988 20244 72268
rect 20076 71932 20244 71988
rect 20076 70756 20132 71932
rect 20076 70700 20244 70756
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19628 69794 19684 69804
rect 20188 70084 20244 70700
rect 20412 70420 20468 72268
rect 20412 70354 20468 70364
rect 19292 69470 19294 69522
rect 19346 69470 19348 69522
rect 19292 69458 19348 69470
rect 19964 69410 20020 69422
rect 19964 69358 19966 69410
rect 20018 69358 20020 69410
rect 19964 69188 20020 69358
rect 19964 69122 20020 69132
rect 19836 69020 20100 69030
rect 19180 68574 19182 68626
rect 19234 68574 19236 68626
rect 19180 68562 19236 68574
rect 19292 68964 19348 68974
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 20188 68964 20244 70028
rect 20524 69636 20580 73838
rect 20748 73890 20804 73902
rect 20748 73838 20750 73890
rect 20802 73838 20804 73890
rect 20636 72436 20692 72446
rect 20636 72342 20692 72380
rect 19292 67058 19348 68908
rect 20188 68898 20244 68908
rect 20300 69580 20580 69636
rect 20076 68180 20132 68190
rect 20076 67954 20132 68124
rect 20076 67902 20078 67954
rect 20130 67902 20132 67954
rect 20076 67890 20132 67902
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 20076 67172 20132 67182
rect 20076 67078 20132 67116
rect 19292 67006 19294 67058
rect 19346 67006 19348 67058
rect 19292 66994 19348 67006
rect 19964 66500 20020 66510
rect 19292 66388 19348 66398
rect 19292 66294 19348 66332
rect 19068 65426 19124 65436
rect 19180 66276 19236 66286
rect 19180 65490 19236 66220
rect 19964 66274 20020 66444
rect 20076 66388 20132 66398
rect 20076 66294 20132 66332
rect 19964 66222 19966 66274
rect 20018 66222 20020 66274
rect 19964 66210 20020 66222
rect 20300 66276 20356 69580
rect 20748 69524 20804 73838
rect 20860 73220 20916 73230
rect 20860 73126 20916 73164
rect 20860 72434 20916 72446
rect 20860 72382 20862 72434
rect 20914 72382 20916 72434
rect 20860 71204 20916 72382
rect 20860 71138 20916 71148
rect 20972 70756 21028 73948
rect 20972 70690 21028 70700
rect 21084 73220 21140 73230
rect 21084 70588 21140 73164
rect 21532 72660 21588 74060
rect 21644 74004 21700 74014
rect 21644 73910 21700 73948
rect 21644 72660 21700 72670
rect 21532 72658 21700 72660
rect 21532 72606 21646 72658
rect 21698 72606 21700 72658
rect 21532 72604 21700 72606
rect 21644 72594 21700 72604
rect 21756 72212 21812 74620
rect 22092 74788 22148 74798
rect 22092 74114 22148 74732
rect 22092 74062 22094 74114
rect 22146 74062 22148 74114
rect 22092 74050 22148 74062
rect 23212 74786 23268 74798
rect 23212 74734 23214 74786
rect 23266 74734 23268 74786
rect 22316 74004 22372 74014
rect 22204 74002 22372 74004
rect 22204 73950 22318 74002
rect 22370 73950 22372 74002
rect 22204 73948 22372 73950
rect 21868 73892 21924 73902
rect 21868 73798 21924 73836
rect 21756 72146 21812 72156
rect 20300 66210 20356 66220
rect 20412 69468 20804 69524
rect 20860 70532 21140 70588
rect 21644 71090 21700 71102
rect 21644 71038 21646 71090
rect 21698 71038 21700 71090
rect 21644 70644 21700 71038
rect 21644 70578 21700 70588
rect 20300 66052 20356 66062
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 20188 65828 20244 65838
rect 19180 65438 19182 65490
rect 19234 65438 19236 65490
rect 19180 65426 19236 65438
rect 19628 65716 19684 65726
rect 19180 65156 19236 65166
rect 18956 64876 19124 64932
rect 18956 64706 19012 64718
rect 18956 64654 18958 64706
rect 19010 64654 19012 64706
rect 18956 64148 19012 64654
rect 18956 64082 19012 64092
rect 18844 63970 18900 63980
rect 19068 64034 19124 64876
rect 19180 64146 19236 65100
rect 19180 64094 19182 64146
rect 19234 64094 19236 64146
rect 19180 64082 19236 64094
rect 19628 64036 19684 65660
rect 20188 65602 20244 65772
rect 20188 65550 20190 65602
rect 20242 65550 20244 65602
rect 20188 65538 20244 65550
rect 20300 65602 20356 65996
rect 20300 65550 20302 65602
rect 20354 65550 20356 65602
rect 19740 65266 19796 65278
rect 19964 65268 20020 65278
rect 19740 65214 19742 65266
rect 19794 65214 19796 65266
rect 19740 64820 19796 65214
rect 19740 64754 19796 64764
rect 19852 65266 20020 65268
rect 19852 65214 19966 65266
rect 20018 65214 20020 65266
rect 19852 65212 20020 65214
rect 19852 64706 19908 65212
rect 19964 65202 20020 65212
rect 19852 64654 19854 64706
rect 19906 64654 19908 64706
rect 19852 64484 19908 64654
rect 20188 64708 20244 64718
rect 20300 64708 20356 65550
rect 20188 64706 20356 64708
rect 20188 64654 20190 64706
rect 20242 64654 20356 64706
rect 20188 64652 20356 64654
rect 20188 64642 20244 64652
rect 19852 64418 19908 64428
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19068 63982 19070 64034
rect 19122 63982 19124 64034
rect 18172 62078 18174 62130
rect 18226 62078 18228 62130
rect 18060 61348 18116 61358
rect 18172 61348 18228 62078
rect 17612 60114 17836 60116
rect 17612 60062 17614 60114
rect 17666 60062 17836 60114
rect 17612 60060 17836 60062
rect 17612 60050 17668 60060
rect 17836 59984 17892 60060
rect 17948 61346 18172 61348
rect 17948 61294 18062 61346
rect 18114 61294 18172 61346
rect 17948 61292 18172 61294
rect 17724 59780 17780 59790
rect 17724 59442 17780 59724
rect 17724 59390 17726 59442
rect 17778 59390 17780 59442
rect 17724 59378 17780 59390
rect 17724 58772 17780 58782
rect 17724 58546 17780 58716
rect 17724 58494 17726 58546
rect 17778 58494 17780 58546
rect 17724 58482 17780 58494
rect 17500 58370 17556 58380
rect 16828 55234 16884 55244
rect 17948 50428 18004 61292
rect 18060 61282 18116 61292
rect 18172 61216 18228 61292
rect 18508 62130 18564 62142
rect 18508 62078 18510 62130
rect 18562 62078 18564 62130
rect 18284 61012 18340 61022
rect 18284 60918 18340 60956
rect 18508 60340 18564 62078
rect 18620 62132 18788 62188
rect 18956 63700 19012 63710
rect 18844 62132 18900 62142
rect 18620 60676 18676 62132
rect 18732 62020 18788 62030
rect 18732 61346 18788 61964
rect 18732 61294 18734 61346
rect 18786 61294 18788 61346
rect 18732 60900 18788 61294
rect 18844 61236 18900 62076
rect 18844 61170 18900 61180
rect 18732 60844 18900 60900
rect 18732 60676 18788 60686
rect 18620 60674 18788 60676
rect 18620 60622 18734 60674
rect 18786 60622 18788 60674
rect 18620 60620 18788 60622
rect 18732 60562 18788 60620
rect 18732 60510 18734 60562
rect 18786 60510 18788 60562
rect 18732 60498 18788 60510
rect 18508 60284 18676 60340
rect 18508 60116 18564 60126
rect 18284 60004 18340 60014
rect 18284 59910 18340 59948
rect 18508 59442 18564 60060
rect 18508 59390 18510 59442
rect 18562 59390 18564 59442
rect 18508 59378 18564 59390
rect 18060 59220 18116 59230
rect 18060 58548 18116 59164
rect 18172 59106 18228 59118
rect 18172 59054 18174 59106
rect 18226 59054 18228 59106
rect 18172 58996 18228 59054
rect 18172 58930 18228 58940
rect 18172 58548 18228 58558
rect 18060 58546 18228 58548
rect 18060 58494 18174 58546
rect 18226 58494 18228 58546
rect 18060 58492 18228 58494
rect 18172 58482 18228 58492
rect 18620 56644 18676 60284
rect 18844 59332 18900 60844
rect 18956 59892 19012 63644
rect 19068 61012 19124 63982
rect 19404 64034 19684 64036
rect 19404 63982 19630 64034
rect 19682 63982 19684 64034
rect 19404 63980 19684 63982
rect 19292 63924 19348 63934
rect 19292 63830 19348 63868
rect 19180 63812 19236 63822
rect 19180 61346 19236 63756
rect 19292 62244 19348 62254
rect 19292 62150 19348 62188
rect 19180 61294 19182 61346
rect 19234 61294 19236 61346
rect 19180 61124 19236 61294
rect 19180 61058 19236 61068
rect 19068 60946 19124 60956
rect 19180 60788 19236 60798
rect 19404 60788 19460 63980
rect 19628 63970 19684 63980
rect 19740 64148 19796 64158
rect 19740 63362 19796 64092
rect 20300 64148 20356 64158
rect 20300 64054 20356 64092
rect 20188 64036 20244 64046
rect 20188 63942 20244 63980
rect 19740 63310 19742 63362
rect 19794 63310 19796 63362
rect 19740 63298 19796 63310
rect 20300 63924 20356 63934
rect 20412 63924 20468 69468
rect 20860 69412 20916 70532
rect 22204 70420 22260 73948
rect 22316 73938 22372 73948
rect 22764 74004 22820 74014
rect 22764 73910 22820 73948
rect 21868 70364 22260 70420
rect 22428 73890 22484 73902
rect 22428 73838 22430 73890
rect 22482 73838 22484 73890
rect 20748 69356 20916 69412
rect 21308 69860 21364 69870
rect 20524 69300 20580 69310
rect 20748 69300 20804 69356
rect 20972 69300 21028 69310
rect 20524 69206 20580 69244
rect 20636 69298 20804 69300
rect 20636 69246 20750 69298
rect 20802 69246 20804 69298
rect 20636 69244 20804 69246
rect 20636 66052 20692 69244
rect 20748 69234 20804 69244
rect 20860 69244 20972 69300
rect 20860 69242 20916 69244
rect 20860 69190 20862 69242
rect 20914 69190 20916 69242
rect 20972 69234 21028 69244
rect 21308 69300 21364 69804
rect 20860 69178 20916 69190
rect 20748 69076 20804 69086
rect 20748 67842 20804 69020
rect 21196 69076 21252 69086
rect 21196 68738 21252 69020
rect 21196 68686 21198 68738
rect 21250 68686 21252 68738
rect 21196 68674 21252 68686
rect 20748 67790 20750 67842
rect 20802 67790 20804 67842
rect 20748 67778 20804 67790
rect 21196 68180 21252 68190
rect 20860 67508 20916 67518
rect 20860 66948 20916 67452
rect 20636 65986 20692 65996
rect 20748 66612 20804 66622
rect 20524 65268 20580 65278
rect 20524 65174 20580 65212
rect 20524 64820 20580 64830
rect 20524 64146 20580 64764
rect 20524 64094 20526 64146
rect 20578 64094 20580 64146
rect 20524 64082 20580 64094
rect 20412 63868 20580 63924
rect 19628 63026 19684 63038
rect 19628 62974 19630 63026
rect 19682 62974 19684 63026
rect 19180 60786 19460 60788
rect 19180 60734 19182 60786
rect 19234 60734 19460 60786
rect 19180 60732 19460 60734
rect 19516 62356 19572 62366
rect 19180 60722 19236 60732
rect 19404 60562 19460 60574
rect 19404 60510 19406 60562
rect 19458 60510 19460 60562
rect 19180 60452 19236 60462
rect 19068 59892 19124 59902
rect 18956 59836 19068 59892
rect 19068 59798 19124 59836
rect 18844 59266 18900 59276
rect 18956 59106 19012 59118
rect 18956 59054 18958 59106
rect 19010 59054 19012 59106
rect 18956 58548 19012 59054
rect 18956 58482 19012 58492
rect 19180 57988 19236 60396
rect 19404 58660 19460 60510
rect 19516 60114 19572 62300
rect 19628 62244 19684 62974
rect 19740 63028 19796 63038
rect 19740 62934 19796 62972
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19740 62580 19796 62590
rect 19740 62486 19796 62524
rect 20188 62580 20244 62590
rect 20300 62580 20356 63868
rect 20188 62578 20356 62580
rect 20188 62526 20190 62578
rect 20242 62526 20356 62578
rect 20188 62524 20356 62526
rect 20412 63252 20468 63262
rect 19628 62178 19684 62188
rect 19740 61572 19796 61582
rect 19740 61478 19796 61516
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19740 61012 19796 61022
rect 20188 61012 20244 62524
rect 20412 61908 20468 63196
rect 20412 61842 20468 61852
rect 20300 61348 20356 61358
rect 20300 61254 20356 61292
rect 20188 60956 20468 61012
rect 19740 60918 19796 60956
rect 20188 60676 20244 60686
rect 20188 60582 20244 60620
rect 19516 60062 19518 60114
rect 19570 60062 19572 60114
rect 19516 60050 19572 60062
rect 20412 60114 20468 60956
rect 20524 60228 20580 63868
rect 20636 63700 20692 63710
rect 20636 62578 20692 63644
rect 20636 62526 20638 62578
rect 20690 62526 20692 62578
rect 20636 62514 20692 62526
rect 20748 62188 20804 66556
rect 20860 66386 20916 66892
rect 20860 66334 20862 66386
rect 20914 66334 20916 66386
rect 20860 65716 20916 66334
rect 20860 65650 20916 65660
rect 20972 65604 21028 65614
rect 20860 64482 20916 64494
rect 20860 64430 20862 64482
rect 20914 64430 20916 64482
rect 20860 64148 20916 64430
rect 20860 64082 20916 64092
rect 20860 62916 20916 62926
rect 20860 62692 20916 62860
rect 20860 62356 20916 62636
rect 20860 62290 20916 62300
rect 20972 62188 21028 65548
rect 21196 64596 21252 68124
rect 21196 64530 21252 64540
rect 21308 65602 21364 69244
rect 21756 69186 21812 69198
rect 21756 69134 21758 69186
rect 21810 69134 21812 69186
rect 21756 68852 21812 69134
rect 21756 68786 21812 68796
rect 21868 68404 21924 70364
rect 22428 70308 22484 73838
rect 22988 73220 23044 73230
rect 22988 73126 23044 73164
rect 21868 68338 21924 68348
rect 21980 70252 22484 70308
rect 22652 71316 22708 71326
rect 21308 65550 21310 65602
rect 21362 65550 21364 65602
rect 21308 64036 21364 65550
rect 21308 63970 21364 63980
rect 21420 67844 21476 67854
rect 21420 63924 21476 67788
rect 21756 67844 21812 67854
rect 21756 67750 21812 67788
rect 21644 67730 21700 67742
rect 21644 67678 21646 67730
rect 21698 67678 21700 67730
rect 21644 67620 21700 67678
rect 21644 67564 21924 67620
rect 21644 67396 21700 67406
rect 21532 67284 21588 67294
rect 21532 65714 21588 67228
rect 21532 65662 21534 65714
rect 21586 65662 21588 65714
rect 21532 64932 21588 65662
rect 21644 65714 21700 67340
rect 21868 66500 21924 67564
rect 21868 66434 21924 66444
rect 21644 65662 21646 65714
rect 21698 65662 21700 65714
rect 21644 65650 21700 65662
rect 21756 66052 21812 66062
rect 21756 65714 21812 65996
rect 21756 65662 21758 65714
rect 21810 65662 21812 65714
rect 21756 65650 21812 65662
rect 21868 65940 21924 65950
rect 21868 65714 21924 65884
rect 21868 65662 21870 65714
rect 21922 65662 21924 65714
rect 21868 65604 21924 65662
rect 21868 65538 21924 65548
rect 21980 65380 22036 70252
rect 22428 70082 22484 70094
rect 22428 70030 22430 70082
rect 22482 70030 22484 70082
rect 22428 69524 22484 70030
rect 22428 69458 22484 69468
rect 22540 69748 22596 69758
rect 22204 69410 22260 69422
rect 22204 69358 22206 69410
rect 22258 69358 22260 69410
rect 22204 69188 22260 69358
rect 22204 69122 22260 69132
rect 22092 67842 22148 67854
rect 22092 67790 22094 67842
rect 22146 67790 22148 67842
rect 22092 67172 22148 67790
rect 22092 67116 22484 67172
rect 22092 67060 22148 67116
rect 22092 66994 22148 67004
rect 22204 66948 22260 66958
rect 22204 66946 22372 66948
rect 22204 66894 22206 66946
rect 22258 66894 22372 66946
rect 22204 66892 22372 66894
rect 22204 66882 22260 66892
rect 21532 64866 21588 64876
rect 21868 65324 22036 65380
rect 22092 66388 22148 66398
rect 21532 63924 21588 63934
rect 21420 63922 21588 63924
rect 21420 63870 21534 63922
rect 21586 63870 21588 63922
rect 21420 63868 21588 63870
rect 21308 63810 21364 63822
rect 21308 63758 21310 63810
rect 21362 63758 21364 63810
rect 21308 63700 21364 63758
rect 21308 63634 21364 63644
rect 21532 62916 21588 63868
rect 21532 62850 21588 62860
rect 21756 63252 21812 63262
rect 21756 63138 21812 63196
rect 21756 63086 21758 63138
rect 21810 63086 21812 63138
rect 21756 62916 21812 63086
rect 21868 63140 21924 65324
rect 22092 64818 22148 66332
rect 22092 64766 22094 64818
rect 22146 64766 22148 64818
rect 22092 64754 22148 64766
rect 22204 66274 22260 66286
rect 22204 66222 22206 66274
rect 22258 66222 22260 66274
rect 22092 64596 22148 64606
rect 21980 64482 22036 64494
rect 21980 64430 21982 64482
rect 22034 64430 22036 64482
rect 21980 63364 22036 64430
rect 21980 63298 22036 63308
rect 22092 63140 22148 64540
rect 22204 64482 22260 66222
rect 22204 64430 22206 64482
rect 22258 64430 22260 64482
rect 22204 64148 22260 64430
rect 22316 64148 22372 66892
rect 22428 64820 22484 67116
rect 22540 65940 22596 69692
rect 22652 67170 22708 71260
rect 22876 70644 22932 70654
rect 22652 67118 22654 67170
rect 22706 67118 22708 67170
rect 22652 67060 22708 67118
rect 22652 66994 22708 67004
rect 22764 70196 22820 70206
rect 22764 66612 22820 70140
rect 22764 66546 22820 66556
rect 22540 65874 22596 65884
rect 22652 66388 22708 66398
rect 22540 65604 22596 65614
rect 22652 65604 22708 66332
rect 22876 66386 22932 70588
rect 23100 70194 23156 70206
rect 23100 70142 23102 70194
rect 23154 70142 23156 70194
rect 22876 66334 22878 66386
rect 22930 66334 22932 66386
rect 22876 66322 22932 66334
rect 22988 69636 23044 69646
rect 22988 69522 23044 69580
rect 22988 69470 22990 69522
rect 23042 69470 23044 69522
rect 22764 66274 22820 66286
rect 22764 66222 22766 66274
rect 22818 66222 22820 66274
rect 22764 66052 22820 66222
rect 22764 65986 22820 65996
rect 22652 65548 22820 65604
rect 22540 65510 22596 65548
rect 22764 65490 22820 65548
rect 22764 65438 22766 65490
rect 22818 65438 22820 65490
rect 22764 65426 22820 65438
rect 22428 64754 22484 64764
rect 22988 64596 23044 69470
rect 23100 69188 23156 70142
rect 23212 70196 23268 74734
rect 23772 74564 23828 74574
rect 23436 74114 23492 74126
rect 23436 74062 23438 74114
rect 23490 74062 23492 74114
rect 23436 72548 23492 74062
rect 23772 73948 23828 74508
rect 24220 74116 24276 74846
rect 24220 74050 24276 74060
rect 24444 74898 24500 74910
rect 24444 74846 24446 74898
rect 24498 74846 24500 74898
rect 24108 74002 24164 74014
rect 24108 73950 24110 74002
rect 24162 73950 24164 74002
rect 23772 73892 23940 73948
rect 23436 72482 23492 72492
rect 23660 73330 23716 73342
rect 23660 73278 23662 73330
rect 23714 73278 23716 73330
rect 23212 70130 23268 70140
rect 23548 70756 23604 70766
rect 23100 69122 23156 69132
rect 23548 67954 23604 70700
rect 23660 70644 23716 73278
rect 23772 72660 23828 72670
rect 23772 72566 23828 72604
rect 23772 71092 23828 71102
rect 23772 70998 23828 71036
rect 23884 70868 23940 73892
rect 23996 73556 24052 73566
rect 24108 73556 24164 73950
rect 23996 73554 24164 73556
rect 23996 73502 23998 73554
rect 24050 73502 24164 73554
rect 23996 73500 24164 73502
rect 23996 73490 24052 73500
rect 24444 73444 24500 74846
rect 24556 73948 24612 78428
rect 24668 75124 24724 79200
rect 27916 78708 27972 78718
rect 25116 78036 25172 78046
rect 24668 75058 24724 75068
rect 24892 75796 24948 75806
rect 24892 75010 24948 75740
rect 25116 75794 25172 77980
rect 27804 77812 27860 77822
rect 27692 77588 27748 77598
rect 27468 77476 27524 77486
rect 27468 76578 27524 77420
rect 27468 76526 27470 76578
rect 27522 76526 27524 76578
rect 27468 76514 27524 76526
rect 25116 75742 25118 75794
rect 25170 75742 25172 75794
rect 25116 75730 25172 75742
rect 25340 76354 25396 76366
rect 25340 76302 25342 76354
rect 25394 76302 25396 76354
rect 24892 74958 24894 75010
rect 24946 74958 24948 75010
rect 24892 74946 24948 74958
rect 24668 74900 24724 74910
rect 24668 74806 24724 74844
rect 24780 74676 24836 74686
rect 24780 74674 25060 74676
rect 24780 74622 24782 74674
rect 24834 74622 25060 74674
rect 24780 74620 25060 74622
rect 24780 74610 24836 74620
rect 24556 73892 24948 73948
rect 24444 73378 24500 73388
rect 24780 73780 24836 73790
rect 23996 73330 24052 73342
rect 23996 73278 23998 73330
rect 24050 73278 24052 73330
rect 23996 72436 24052 73278
rect 24332 73330 24388 73342
rect 24332 73278 24334 73330
rect 24386 73278 24388 73330
rect 24332 72772 24388 73278
rect 24332 72706 24388 72716
rect 23996 72370 24052 72380
rect 24444 72548 24500 72558
rect 24220 71650 24276 71662
rect 24220 71598 24222 71650
rect 24274 71598 24276 71650
rect 24220 70980 24276 71598
rect 24444 70980 24500 72492
rect 24780 71764 24836 73724
rect 24892 73218 24948 73892
rect 24892 73166 24894 73218
rect 24946 73166 24948 73218
rect 24892 71988 24948 73166
rect 24892 71922 24948 71932
rect 24892 71764 24948 71774
rect 24780 71762 24948 71764
rect 24780 71710 24894 71762
rect 24946 71710 24948 71762
rect 24780 71708 24948 71710
rect 24556 70980 24612 70990
rect 24220 70978 24724 70980
rect 24220 70926 24558 70978
rect 24610 70926 24724 70978
rect 24220 70924 24724 70926
rect 24556 70914 24612 70924
rect 23660 70578 23716 70588
rect 23772 70812 24164 70868
rect 23548 67902 23550 67954
rect 23602 67902 23604 67954
rect 23548 67890 23604 67902
rect 23436 67844 23492 67854
rect 23436 67750 23492 67788
rect 23660 67844 23716 67854
rect 23772 67844 23828 70812
rect 23884 70644 23940 70654
rect 23884 70418 23940 70588
rect 23884 70366 23886 70418
rect 23938 70366 23940 70418
rect 23884 70354 23940 70366
rect 24108 70418 24164 70812
rect 24332 70756 24388 70766
rect 24332 70588 24388 70700
rect 24332 70532 24612 70588
rect 24108 70366 24110 70418
rect 24162 70366 24164 70418
rect 24108 70354 24164 70366
rect 24332 70196 24388 70206
rect 24332 70102 24388 70140
rect 24220 70082 24276 70094
rect 24220 70030 24222 70082
rect 24274 70030 24276 70082
rect 24108 68404 24164 68414
rect 23660 67842 23828 67844
rect 23660 67790 23662 67842
rect 23714 67790 23828 67842
rect 23660 67788 23828 67790
rect 23660 67778 23716 67788
rect 23212 67730 23268 67742
rect 23212 67678 23214 67730
rect 23266 67678 23268 67730
rect 23212 67620 23268 67678
rect 23212 67554 23268 67564
rect 23548 66500 23604 66510
rect 23436 66388 23492 66398
rect 23212 66386 23492 66388
rect 23212 66334 23438 66386
rect 23490 66334 23492 66386
rect 23212 66332 23492 66334
rect 23100 64820 23156 64830
rect 23100 64726 23156 64764
rect 22988 64540 23156 64596
rect 22428 64484 22484 64494
rect 22428 64390 22484 64428
rect 22988 64260 23044 64270
rect 22764 64148 22820 64158
rect 22316 64146 22820 64148
rect 22316 64094 22766 64146
rect 22818 64094 22820 64146
rect 22316 64092 22820 64094
rect 22204 64082 22260 64092
rect 22764 64082 22820 64092
rect 22204 63924 22260 63934
rect 22204 63830 22260 63868
rect 22988 63924 23044 64204
rect 22316 63588 22372 63598
rect 22092 63084 22260 63140
rect 21868 63008 21924 63084
rect 21756 62850 21812 62860
rect 21980 62914 22036 62926
rect 21980 62862 21982 62914
rect 22034 62862 22036 62914
rect 21084 62804 21140 62814
rect 21084 62578 21140 62748
rect 21084 62526 21086 62578
rect 21138 62526 21140 62578
rect 21084 62514 21140 62526
rect 21532 62580 21588 62590
rect 21532 62486 21588 62524
rect 20636 62132 20804 62188
rect 20860 62132 21028 62188
rect 21980 62244 22036 62862
rect 22092 62914 22148 62926
rect 22092 62862 22094 62914
rect 22146 62862 22148 62914
rect 22092 62804 22148 62862
rect 22204 62916 22260 63084
rect 22316 63138 22372 63532
rect 22876 63364 22932 63374
rect 22876 63270 22932 63308
rect 22988 63250 23044 63868
rect 22988 63198 22990 63250
rect 23042 63198 23044 63250
rect 22988 63186 23044 63198
rect 22316 63086 22318 63138
rect 22370 63086 22372 63138
rect 22316 63074 22372 63086
rect 22764 63140 22820 63150
rect 22204 62860 22484 62916
rect 22092 62738 22148 62748
rect 22092 62580 22148 62590
rect 22092 62466 22148 62524
rect 22092 62414 22094 62466
rect 22146 62414 22148 62466
rect 22092 62402 22148 62414
rect 22204 62468 22260 62478
rect 22260 62412 22372 62468
rect 22204 62374 22260 62412
rect 21980 62178 22036 62188
rect 20636 61010 20692 62132
rect 20748 61684 20804 61694
rect 20860 61684 20916 62132
rect 21868 61794 21924 61806
rect 21868 61742 21870 61794
rect 21922 61742 21924 61794
rect 20748 61682 20916 61684
rect 20748 61630 20750 61682
rect 20802 61630 20916 61682
rect 20748 61628 20916 61630
rect 21756 61684 21812 61694
rect 20748 61618 20804 61628
rect 21756 61590 21812 61628
rect 20636 60958 20638 61010
rect 20690 60958 20692 61010
rect 20636 60946 20692 60958
rect 21308 61348 21364 61358
rect 21308 60674 21364 61292
rect 21868 61010 21924 61742
rect 21868 60958 21870 61010
rect 21922 60958 21924 61010
rect 21868 60946 21924 60958
rect 22204 61796 22260 61806
rect 22204 61682 22260 61740
rect 22204 61630 22206 61682
rect 22258 61630 22260 61682
rect 21308 60622 21310 60674
rect 21362 60622 21364 60674
rect 20524 60162 20580 60172
rect 20860 60452 20916 60462
rect 20412 60062 20414 60114
rect 20466 60062 20468 60114
rect 20412 60050 20468 60062
rect 20860 60114 20916 60396
rect 20860 60062 20862 60114
rect 20914 60062 20916 60114
rect 19852 59780 19908 59790
rect 19516 59778 19908 59780
rect 19516 59726 19854 59778
rect 19906 59726 19908 59778
rect 19516 59724 19908 59726
rect 19516 58996 19572 59724
rect 19852 59714 19908 59724
rect 20860 59780 20916 60062
rect 20860 59714 20916 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 21308 59444 21364 60622
rect 22204 60452 22260 61630
rect 22316 61012 22372 62412
rect 22428 61794 22484 62860
rect 22428 61742 22430 61794
rect 22482 61742 22484 61794
rect 22428 61730 22484 61742
rect 22540 62804 22596 62814
rect 22540 61012 22596 62748
rect 22764 62578 22820 63084
rect 22764 62526 22766 62578
rect 22818 62526 22820 62578
rect 22764 62514 22820 62526
rect 22652 62244 22708 62254
rect 23100 62188 23156 64540
rect 23212 63476 23268 66332
rect 23436 66322 23492 66332
rect 23436 66052 23492 66062
rect 23436 65490 23492 65996
rect 23548 65602 23604 66444
rect 23548 65550 23550 65602
rect 23602 65550 23604 65602
rect 23548 65538 23604 65550
rect 23436 65438 23438 65490
rect 23490 65438 23492 65490
rect 23324 64820 23380 64830
rect 23324 64036 23380 64764
rect 23436 64260 23492 65438
rect 23772 65380 23828 67788
rect 23884 67844 23940 67854
rect 23884 67750 23940 67788
rect 24108 67508 24164 68348
rect 23772 65314 23828 65324
rect 23884 67058 23940 67070
rect 23884 67006 23886 67058
rect 23938 67006 23940 67058
rect 23884 65602 23940 67006
rect 23996 66948 24052 66958
rect 23996 66854 24052 66892
rect 23884 65550 23886 65602
rect 23938 65550 23940 65602
rect 23884 65044 23940 65550
rect 23884 64978 23940 64988
rect 23436 64194 23492 64204
rect 23548 64932 23604 64942
rect 23436 64036 23492 64046
rect 23324 64034 23436 64036
rect 23324 63982 23326 64034
rect 23378 63982 23436 64034
rect 23324 63980 23436 63982
rect 23324 63970 23380 63980
rect 23212 63410 23268 63420
rect 23324 63588 23380 63598
rect 23324 62578 23380 63532
rect 23324 62526 23326 62578
rect 23378 62526 23380 62578
rect 23324 62514 23380 62526
rect 23436 62356 23492 63980
rect 22652 61348 22708 62188
rect 22652 61254 22708 61292
rect 22764 62132 23156 62188
rect 23212 62300 23492 62356
rect 22652 61012 22708 61022
rect 22540 61010 22708 61012
rect 22540 60958 22654 61010
rect 22706 60958 22708 61010
rect 22540 60956 22708 60958
rect 22316 60880 22372 60956
rect 22652 60946 22708 60956
rect 22764 60788 22820 62132
rect 23100 61346 23156 61358
rect 23100 61294 23102 61346
rect 23154 61294 23156 61346
rect 23100 61236 23156 61294
rect 23100 61170 23156 61180
rect 22204 60386 22260 60396
rect 22428 60732 22820 60788
rect 22428 60228 22484 60732
rect 23212 60676 23268 62300
rect 23548 62188 23604 64876
rect 23772 64932 23828 64942
rect 23772 64706 23828 64876
rect 23996 64820 24052 64830
rect 23996 64726 24052 64764
rect 23772 64654 23774 64706
rect 23826 64654 23828 64706
rect 23772 64642 23828 64654
rect 23884 64708 23940 64718
rect 23884 63924 23940 64652
rect 24108 64706 24164 67452
rect 24220 67284 24276 70030
rect 24220 67218 24276 67228
rect 24332 69636 24388 69646
rect 24332 67170 24388 69580
rect 24444 68516 24500 68526
rect 24444 67956 24500 68460
rect 24444 67842 24500 67900
rect 24444 67790 24446 67842
rect 24498 67790 24500 67842
rect 24444 67778 24500 67790
rect 24556 67620 24612 70532
rect 24332 67118 24334 67170
rect 24386 67118 24388 67170
rect 24332 67106 24388 67118
rect 24444 67508 24500 67518
rect 24444 66388 24500 67452
rect 24332 66332 24500 66388
rect 24220 65492 24276 65502
rect 24220 65398 24276 65436
rect 24108 64654 24110 64706
rect 24162 64654 24164 64706
rect 24108 64642 24164 64654
rect 24332 64708 24388 66332
rect 24444 65268 24500 65278
rect 24444 65174 24500 65212
rect 24332 64706 24500 64708
rect 24332 64654 24334 64706
rect 24386 64654 24500 64706
rect 24332 64652 24500 64654
rect 24332 64642 24388 64652
rect 24332 64484 24388 64494
rect 24108 64148 24164 64158
rect 24108 64054 24164 64092
rect 23772 63868 23884 63924
rect 23660 63700 23716 63710
rect 23660 63252 23716 63644
rect 23660 63120 23716 63196
rect 23436 62132 23604 62188
rect 23660 62692 23716 62702
rect 23436 61236 23492 62132
rect 23548 62020 23604 62030
rect 23548 61682 23604 61964
rect 23548 61630 23550 61682
rect 23602 61630 23604 61682
rect 23548 61618 23604 61630
rect 23436 61170 23492 61180
rect 23548 61012 23604 61022
rect 23660 61012 23716 62636
rect 23772 62578 23828 63868
rect 23884 63858 23940 63868
rect 23884 63698 23940 63710
rect 23884 63646 23886 63698
rect 23938 63646 23940 63698
rect 23884 63364 23940 63646
rect 24220 63700 24276 63710
rect 24220 63606 24276 63644
rect 23884 63298 23940 63308
rect 24108 63476 24164 63486
rect 23772 62526 23774 62578
rect 23826 62526 23828 62578
rect 23772 62514 23828 62526
rect 23548 61010 23716 61012
rect 23548 60958 23550 61010
rect 23602 60958 23716 61010
rect 23548 60956 23716 60958
rect 23772 62020 23828 62030
rect 23772 61684 23828 61964
rect 23548 60946 23604 60956
rect 23212 60582 23268 60620
rect 21980 60172 22484 60228
rect 21980 60114 22036 60172
rect 21980 60062 21982 60114
rect 22034 60062 22036 60114
rect 21980 60050 22036 60062
rect 23212 60116 23268 60126
rect 23212 60022 23268 60060
rect 23660 60116 23716 60126
rect 23772 60116 23828 61628
rect 24108 61010 24164 63420
rect 24332 63364 24388 64428
rect 24220 63252 24276 63262
rect 24332 63232 24388 63308
rect 24220 63138 24276 63196
rect 24220 63086 24222 63138
rect 24274 63086 24276 63138
rect 24220 63074 24276 63086
rect 24332 62916 24388 62926
rect 24220 62914 24388 62916
rect 24220 62862 24334 62914
rect 24386 62862 24388 62914
rect 24220 62860 24388 62862
rect 24220 62692 24276 62860
rect 24332 62850 24388 62860
rect 24220 62626 24276 62636
rect 24332 62580 24388 62590
rect 24444 62580 24500 64652
rect 24556 63476 24612 67564
rect 24556 63410 24612 63420
rect 24668 63140 24724 70924
rect 24892 70308 24948 71708
rect 24780 70252 24892 70308
rect 24780 68404 24836 70252
rect 24892 70242 24948 70252
rect 24892 70082 24948 70094
rect 24892 70030 24894 70082
rect 24946 70030 24948 70082
rect 24892 69972 24948 70030
rect 24892 68850 24948 69916
rect 24892 68798 24894 68850
rect 24946 68798 24948 68850
rect 24892 68786 24948 68798
rect 24780 68338 24836 68348
rect 24780 67956 24836 67966
rect 24780 67842 24836 67900
rect 24780 67790 24782 67842
rect 24834 67790 24836 67842
rect 24780 67778 24836 67790
rect 25004 67172 25060 74620
rect 25116 73108 25172 73118
rect 25116 72658 25172 73052
rect 25116 72606 25118 72658
rect 25170 72606 25172 72658
rect 25116 72594 25172 72606
rect 25340 71428 25396 76302
rect 27132 76132 27188 76142
rect 25788 75460 25844 75470
rect 25788 75366 25844 75404
rect 27020 75012 27076 75022
rect 25676 74788 25732 74798
rect 25676 74694 25732 74732
rect 25340 71362 25396 71372
rect 25564 74676 25620 74686
rect 25228 71204 25284 71214
rect 25228 71110 25284 71148
rect 25564 70978 25620 74620
rect 26348 74226 26404 74238
rect 26348 74174 26350 74226
rect 26402 74174 26404 74226
rect 26348 73668 26404 74174
rect 27020 74226 27076 74956
rect 27020 74174 27022 74226
rect 27074 74174 27076 74226
rect 26348 73602 26404 73612
rect 26684 73668 26740 73678
rect 26124 73556 26180 73566
rect 25676 73220 25732 73230
rect 25676 73126 25732 73164
rect 25788 72324 25844 72334
rect 25788 72230 25844 72268
rect 25676 71764 25732 71774
rect 25676 71670 25732 71708
rect 25900 71762 25956 71774
rect 25900 71710 25902 71762
rect 25954 71710 25956 71762
rect 25564 70926 25566 70978
rect 25618 70926 25620 70978
rect 25564 70914 25620 70926
rect 25788 71650 25844 71662
rect 25788 71598 25790 71650
rect 25842 71598 25844 71650
rect 25116 70866 25172 70878
rect 25116 70814 25118 70866
rect 25170 70814 25172 70866
rect 25116 70532 25172 70814
rect 25452 70868 25508 70878
rect 25452 70774 25508 70812
rect 25116 70196 25172 70476
rect 25788 70420 25844 71598
rect 25116 70130 25172 70140
rect 25452 70364 25844 70420
rect 25116 69522 25172 69534
rect 25116 69470 25118 69522
rect 25170 69470 25172 69522
rect 25116 69300 25172 69470
rect 25116 69234 25172 69244
rect 24780 67116 25060 67172
rect 25340 69188 25396 69198
rect 25340 67842 25396 69132
rect 25452 68180 25508 70364
rect 25900 70308 25956 71710
rect 26124 71202 26180 73500
rect 26572 72212 26628 72222
rect 26348 71876 26404 71886
rect 26348 71762 26404 71820
rect 26348 71710 26350 71762
rect 26402 71710 26404 71762
rect 26348 71698 26404 71710
rect 26124 71150 26126 71202
rect 26178 71150 26180 71202
rect 26124 71138 26180 71150
rect 26236 71540 26292 71550
rect 26236 71202 26292 71484
rect 26572 71540 26628 72156
rect 26572 71474 26628 71484
rect 26236 71150 26238 71202
rect 26290 71150 26292 71202
rect 26236 71138 26292 71150
rect 26460 70866 26516 70878
rect 26460 70814 26462 70866
rect 26514 70814 26516 70866
rect 25452 68114 25508 68124
rect 25564 70252 25956 70308
rect 26012 70756 26068 70766
rect 25564 68068 25620 70252
rect 25676 70084 25732 70094
rect 25676 69990 25732 70028
rect 26012 69972 26068 70700
rect 25788 69916 26068 69972
rect 26460 69972 26516 70814
rect 25788 69524 25844 69916
rect 25676 69468 25844 69524
rect 26012 69748 26068 69758
rect 25676 68852 25732 69468
rect 25788 69186 25844 69198
rect 25788 69134 25790 69186
rect 25842 69134 25844 69186
rect 25788 68852 25844 69134
rect 26012 69186 26068 69692
rect 26460 69524 26516 69916
rect 26460 69458 26516 69468
rect 26572 70084 26628 70094
rect 26124 69412 26180 69422
rect 26124 69318 26180 69356
rect 26012 69134 26014 69186
rect 26066 69134 26068 69186
rect 26012 69076 26068 69134
rect 26236 69188 26292 69198
rect 26236 69186 26516 69188
rect 26236 69134 26238 69186
rect 26290 69134 26516 69186
rect 26236 69132 26516 69134
rect 26236 69122 26292 69132
rect 26012 69010 26068 69020
rect 26124 68964 26180 68974
rect 26012 68852 26068 68862
rect 25788 68850 26068 68852
rect 25788 68798 26014 68850
rect 26066 68798 26068 68850
rect 25788 68796 26068 68798
rect 25676 68738 25732 68796
rect 26012 68786 26068 68796
rect 26124 68850 26180 68908
rect 26124 68798 26126 68850
rect 26178 68798 26180 68850
rect 26124 68786 26180 68798
rect 26348 68852 26404 68862
rect 25676 68686 25678 68738
rect 25730 68686 25732 68738
rect 25676 68674 25732 68686
rect 25900 68626 25956 68638
rect 25900 68574 25902 68626
rect 25954 68574 25956 68626
rect 25900 68404 25956 68574
rect 25900 68338 25956 68348
rect 26012 68628 26068 68638
rect 25564 68002 25620 68012
rect 26012 67954 26068 68572
rect 26012 67902 26014 67954
rect 26066 67902 26068 67954
rect 26012 67890 26068 67902
rect 26236 68628 26292 68638
rect 25340 67790 25342 67842
rect 25394 67790 25396 67842
rect 24780 63588 24836 67116
rect 24892 66946 24948 66958
rect 24892 66894 24894 66946
rect 24946 66894 24948 66946
rect 24892 65940 24948 66894
rect 25340 66612 25396 67790
rect 25788 67508 25844 67518
rect 26236 67508 26292 68572
rect 25676 67058 25732 67070
rect 25676 67006 25678 67058
rect 25730 67006 25732 67058
rect 25340 66546 25396 66556
rect 25452 66948 25508 66958
rect 24892 65714 24948 65884
rect 25452 66276 25508 66892
rect 24892 65662 24894 65714
rect 24946 65662 24948 65714
rect 24892 65604 24948 65662
rect 24892 65538 24948 65548
rect 25116 65716 25172 65726
rect 24780 63522 24836 63532
rect 24892 65380 24948 65390
rect 24892 64260 24948 65324
rect 25116 65156 25172 65660
rect 25116 65090 25172 65100
rect 25116 64708 25172 64718
rect 24892 64146 24948 64204
rect 24892 64094 24894 64146
rect 24946 64094 24948 64146
rect 24332 62578 24500 62580
rect 24332 62526 24334 62578
rect 24386 62526 24500 62578
rect 24332 62524 24500 62526
rect 24556 63084 24724 63140
rect 24332 62514 24388 62524
rect 24220 61684 24276 61694
rect 24220 61590 24276 61628
rect 24556 61684 24612 63084
rect 24668 62692 24724 62702
rect 24668 62578 24724 62636
rect 24668 62526 24670 62578
rect 24722 62526 24724 62578
rect 24668 62514 24724 62526
rect 24892 62020 24948 64094
rect 25004 64652 25116 64708
rect 25004 63364 25060 64652
rect 25116 64614 25172 64652
rect 25340 64706 25396 64718
rect 25340 64654 25342 64706
rect 25394 64654 25396 64706
rect 25340 64036 25396 64654
rect 25452 64596 25508 66220
rect 25564 66164 25620 66174
rect 25564 66070 25620 66108
rect 25676 64820 25732 67006
rect 25676 64754 25732 64764
rect 25452 64530 25508 64540
rect 25676 64596 25732 64606
rect 25676 64502 25732 64540
rect 25564 64482 25620 64494
rect 25564 64430 25566 64482
rect 25618 64430 25620 64482
rect 25564 64372 25620 64430
rect 25788 64484 25844 67452
rect 25900 67452 26292 67508
rect 25900 64932 25956 67452
rect 26348 67396 26404 68796
rect 26348 67330 26404 67340
rect 26236 67284 26292 67294
rect 26124 67172 26180 67182
rect 26124 67078 26180 67116
rect 26236 67170 26292 67228
rect 26236 67118 26238 67170
rect 26290 67118 26292 67170
rect 26236 67106 26292 67118
rect 26012 67058 26068 67070
rect 26012 67006 26014 67058
rect 26066 67006 26068 67058
rect 26012 66052 26068 67006
rect 26236 66612 26292 66622
rect 26236 66274 26292 66556
rect 26236 66222 26238 66274
rect 26290 66222 26292 66274
rect 26236 66210 26292 66222
rect 26460 66164 26516 69132
rect 26572 68964 26628 70028
rect 26684 69636 26740 73612
rect 26796 71538 26852 71550
rect 26796 71486 26798 71538
rect 26850 71486 26852 71538
rect 26796 70084 26852 71486
rect 26908 71540 26964 71550
rect 26908 71446 26964 71484
rect 27020 71428 27076 74174
rect 27020 71362 27076 71372
rect 27132 74116 27188 76076
rect 27132 71090 27188 74060
rect 27356 73556 27412 73566
rect 27132 71038 27134 71090
rect 27186 71038 27188 71090
rect 27132 71026 27188 71038
rect 27244 73332 27300 73342
rect 27244 71986 27300 73276
rect 27244 71934 27246 71986
rect 27298 71934 27300 71986
rect 27244 70868 27300 71934
rect 27244 70802 27300 70812
rect 26796 70018 26852 70028
rect 26684 69580 26964 69636
rect 26572 68898 26628 68908
rect 26796 69410 26852 69422
rect 26796 69358 26798 69410
rect 26850 69358 26852 69410
rect 26796 68964 26852 69358
rect 26796 68898 26852 68908
rect 26908 68740 26964 69580
rect 27356 69524 27412 73500
rect 27692 71988 27748 77532
rect 27804 75010 27860 77756
rect 27804 74958 27806 75010
rect 27858 74958 27860 75010
rect 27804 74946 27860 74958
rect 27916 77700 27972 78652
rect 27804 73220 27860 73230
rect 27804 73126 27860 73164
rect 27916 72660 27972 77644
rect 28028 77588 28084 77598
rect 28028 75794 28084 77532
rect 28588 77588 28644 79548
rect 28588 77522 28644 77532
rect 28140 76468 28196 76478
rect 28140 76374 28196 76412
rect 28700 76468 28756 76478
rect 28028 75742 28030 75794
rect 28082 75742 28084 75794
rect 28028 75730 28084 75742
rect 28364 75908 28420 75918
rect 28364 75124 28420 75852
rect 28364 74002 28420 75068
rect 28700 75682 28756 76412
rect 28700 75630 28702 75682
rect 28754 75630 28756 75682
rect 28364 73950 28366 74002
rect 28418 73950 28420 74002
rect 28364 73938 28420 73950
rect 28588 74900 28644 74910
rect 28700 74900 28756 75630
rect 28588 74898 28756 74900
rect 28588 74846 28590 74898
rect 28642 74846 28756 74898
rect 28588 74844 28756 74846
rect 28588 73330 28644 74844
rect 28812 73948 28868 79660
rect 29008 79200 29120 80000
rect 33376 79200 33488 80000
rect 37744 79200 37856 80000
rect 42112 79200 42224 80000
rect 46480 79200 46592 80000
rect 50848 79200 50960 80000
rect 55216 79200 55328 80000
rect 59584 79200 59696 80000
rect 63952 79200 64064 80000
rect 68320 79200 68432 80000
rect 72688 79200 72800 80000
rect 77056 79200 77168 80000
rect 29036 75348 29092 79200
rect 31836 76916 31892 76926
rect 31724 76692 31780 76702
rect 30604 76578 30660 76590
rect 30604 76526 30606 76578
rect 30658 76526 30660 76578
rect 29484 76356 29540 76366
rect 29484 76354 29988 76356
rect 29484 76302 29486 76354
rect 29538 76302 29988 76354
rect 29484 76300 29988 76302
rect 29484 76290 29540 76300
rect 29820 75796 29876 75806
rect 29820 75702 29876 75740
rect 29036 75282 29092 75292
rect 29708 74898 29764 74910
rect 29708 74846 29710 74898
rect 29762 74846 29764 74898
rect 28588 73278 28590 73330
rect 28642 73278 28644 73330
rect 28028 72660 28084 72670
rect 27916 72658 28084 72660
rect 27916 72606 28030 72658
rect 28082 72606 28084 72658
rect 27916 72604 28084 72606
rect 28028 72594 28084 72604
rect 28588 72548 28644 73278
rect 28588 72482 28644 72492
rect 28700 73892 28868 73948
rect 29036 74786 29092 74798
rect 29036 74734 29038 74786
rect 29090 74734 29092 74786
rect 29036 73948 29092 74734
rect 29708 73948 29764 74846
rect 28924 73892 28980 73902
rect 29036 73892 29316 73948
rect 28700 72324 28756 73892
rect 28812 73556 28868 73566
rect 28812 73220 28868 73500
rect 28812 73154 28868 73164
rect 28812 72548 28868 72558
rect 28812 72454 28868 72492
rect 28588 72268 28756 72324
rect 28252 72212 28308 72222
rect 27692 71932 27860 71988
rect 27468 71762 27524 71774
rect 27468 71710 27470 71762
rect 27522 71710 27524 71762
rect 27468 71316 27524 71710
rect 27580 71764 27636 71774
rect 27580 71670 27636 71708
rect 27692 71762 27748 71774
rect 27692 71710 27694 71762
rect 27746 71710 27748 71762
rect 27468 71250 27524 71260
rect 27580 70978 27636 70990
rect 27580 70926 27582 70978
rect 27634 70926 27636 70978
rect 27580 70532 27636 70926
rect 27580 69860 27636 70476
rect 27580 69794 27636 69804
rect 27692 70644 27748 71710
rect 27356 69468 27524 69524
rect 27132 69412 27188 69422
rect 27132 69318 27188 69356
rect 26796 68684 26964 68740
rect 27244 69186 27300 69198
rect 27244 69134 27246 69186
rect 27298 69134 27300 69186
rect 26796 67508 26852 68684
rect 27244 68626 27300 69134
rect 27244 68574 27246 68626
rect 27298 68574 27300 68626
rect 27244 68562 27300 68574
rect 27356 69186 27412 69198
rect 27356 69134 27358 69186
rect 27410 69134 27412 69186
rect 26908 68404 26964 68414
rect 26908 68402 27076 68404
rect 26908 68350 26910 68402
rect 26962 68350 27076 68402
rect 26908 68348 27076 68350
rect 26908 68338 26964 68348
rect 26796 67442 26852 67452
rect 26908 67170 26964 67182
rect 26908 67118 26910 67170
rect 26962 67118 26964 67170
rect 26796 67060 26852 67070
rect 26796 66966 26852 67004
rect 26908 66500 26964 67118
rect 26796 66444 26964 66500
rect 26460 66108 26740 66164
rect 26012 65986 26068 65996
rect 26684 65940 26740 66108
rect 26796 66052 26852 66444
rect 27020 66388 27076 68348
rect 27356 67956 27412 69134
rect 27356 67890 27412 67900
rect 27468 68626 27524 69468
rect 27468 68574 27470 68626
rect 27522 68574 27524 68626
rect 27468 67844 27524 68574
rect 27468 67778 27524 67788
rect 27132 67172 27188 67182
rect 27132 67078 27188 67116
rect 27020 66322 27076 66332
rect 27356 66836 27412 66846
rect 27580 66836 27636 66846
rect 26908 66276 26964 66286
rect 26908 66182 26964 66220
rect 27132 66276 27188 66286
rect 27132 66182 27188 66220
rect 26796 65996 26964 66052
rect 26684 65884 26852 65940
rect 26684 65602 26740 65614
rect 26684 65550 26686 65602
rect 26738 65550 26740 65602
rect 26012 65492 26068 65502
rect 26012 65398 26068 65436
rect 26460 65492 26516 65502
rect 26460 65398 26516 65436
rect 25900 64866 25956 64876
rect 26348 65380 26404 65390
rect 26348 65156 26404 65324
rect 26684 65380 26740 65550
rect 26684 65314 26740 65324
rect 26348 64706 26404 65100
rect 26348 64654 26350 64706
rect 26402 64654 26404 64706
rect 26348 64642 26404 64654
rect 26684 64708 26740 64718
rect 26684 64614 26740 64652
rect 25788 64482 25956 64484
rect 25788 64430 25790 64482
rect 25842 64430 25956 64482
rect 25788 64428 25956 64430
rect 25788 64418 25844 64428
rect 25564 64316 25732 64372
rect 25116 63980 25396 64036
rect 25676 64036 25732 64316
rect 25788 64036 25844 64046
rect 25676 63980 25788 64036
rect 25116 63700 25172 63980
rect 25564 63924 25620 63934
rect 25116 63634 25172 63644
rect 25228 63922 25620 63924
rect 25228 63870 25566 63922
rect 25618 63870 25620 63922
rect 25228 63868 25620 63870
rect 25116 63364 25172 63374
rect 25004 63362 25172 63364
rect 25004 63310 25118 63362
rect 25170 63310 25172 63362
rect 25004 63308 25172 63310
rect 25116 63298 25172 63308
rect 25116 63140 25172 63150
rect 25116 63026 25172 63084
rect 25228 63138 25284 63868
rect 25564 63858 25620 63868
rect 25228 63086 25230 63138
rect 25282 63086 25284 63138
rect 25228 63074 25284 63086
rect 25116 62974 25118 63026
rect 25170 62974 25172 63026
rect 25116 62962 25172 62974
rect 25564 62580 25620 62590
rect 25676 62580 25732 63980
rect 25788 63942 25844 63980
rect 25900 64034 25956 64428
rect 25900 63982 25902 64034
rect 25954 63982 25956 64034
rect 25900 63812 25956 63982
rect 26572 64148 26628 64158
rect 26460 63924 26516 63934
rect 26572 63924 26628 64092
rect 26796 64146 26852 65884
rect 26908 65268 26964 65996
rect 27020 66050 27076 66062
rect 27020 65998 27022 66050
rect 27074 65998 27076 66050
rect 27020 65492 27076 65998
rect 27356 65716 27412 66780
rect 27356 65602 27412 65660
rect 27356 65550 27358 65602
rect 27410 65550 27412 65602
rect 27356 65538 27412 65550
rect 27468 66834 27636 66836
rect 27468 66782 27582 66834
rect 27634 66782 27636 66834
rect 27468 66780 27636 66782
rect 27468 65604 27524 66780
rect 27580 66770 27636 66780
rect 27468 65538 27524 65548
rect 27580 66274 27636 66286
rect 27580 66222 27582 66274
rect 27634 66222 27636 66274
rect 27020 65426 27076 65436
rect 27580 65492 27636 66222
rect 27580 65426 27636 65436
rect 27692 65490 27748 70588
rect 27804 70082 27860 71932
rect 27804 70030 27806 70082
rect 27858 70030 27860 70082
rect 27804 68292 27860 70030
rect 28028 70866 28084 70878
rect 28028 70814 28030 70866
rect 28082 70814 28084 70866
rect 28028 69636 28084 70814
rect 28140 69636 28196 69646
rect 28028 69634 28196 69636
rect 28028 69582 28142 69634
rect 28194 69582 28196 69634
rect 28028 69580 28196 69582
rect 28028 69412 28084 69422
rect 28028 69318 28084 69356
rect 27804 68226 27860 68236
rect 28028 68852 28084 68862
rect 28028 67508 28084 68796
rect 28140 68628 28196 69580
rect 28252 68852 28308 72156
rect 28364 71650 28420 71662
rect 28364 71598 28366 71650
rect 28418 71598 28420 71650
rect 28364 69636 28420 71598
rect 28588 71202 28644 72268
rect 28924 72212 28980 73836
rect 29148 73444 29204 73454
rect 29148 73350 29204 73388
rect 29148 73106 29204 73118
rect 29148 73054 29150 73106
rect 29202 73054 29204 73106
rect 29036 72772 29092 72782
rect 29148 72772 29204 73054
rect 29092 72716 29204 72772
rect 29036 72706 29092 72716
rect 29260 72660 29316 73892
rect 29596 73892 29764 73948
rect 29932 74228 29988 76300
rect 30492 75796 30548 75806
rect 30380 74900 30436 74910
rect 29372 73332 29428 73342
rect 29372 73238 29428 73276
rect 28700 72156 28980 72212
rect 28700 71762 28756 72156
rect 28700 71710 28702 71762
rect 28754 71710 28756 71762
rect 28700 71698 28756 71710
rect 28812 71988 28868 71998
rect 28588 71150 28590 71202
rect 28642 71150 28644 71202
rect 28588 71138 28644 71150
rect 28700 71092 28756 71102
rect 28812 71092 28868 71932
rect 28700 71090 28868 71092
rect 28700 71038 28702 71090
rect 28754 71038 28868 71090
rect 28700 71036 28868 71038
rect 28700 71026 28756 71036
rect 28364 69570 28420 69580
rect 28588 70194 28644 70206
rect 28588 70142 28590 70194
rect 28642 70142 28644 70194
rect 28588 69636 28644 70142
rect 28588 69570 28644 69580
rect 28364 69410 28420 69422
rect 28364 69358 28366 69410
rect 28418 69358 28420 69410
rect 28364 69076 28420 69358
rect 28588 69412 28644 69422
rect 28588 69318 28644 69356
rect 28812 69410 28868 69422
rect 28812 69358 28814 69410
rect 28866 69358 28868 69410
rect 28364 69010 28420 69020
rect 28476 69300 28532 69310
rect 28252 68786 28308 68796
rect 28252 68628 28308 68638
rect 28140 68626 28308 68628
rect 28140 68574 28254 68626
rect 28306 68574 28308 68626
rect 28140 68572 28308 68574
rect 28252 68562 28308 68572
rect 28140 67956 28196 67966
rect 28140 67954 28420 67956
rect 28140 67902 28142 67954
rect 28194 67902 28420 67954
rect 28140 67900 28420 67902
rect 28140 67890 28196 67900
rect 27916 67058 27972 67070
rect 27916 67006 27918 67058
rect 27970 67006 27972 67058
rect 27804 66946 27860 66958
rect 27804 66894 27806 66946
rect 27858 66894 27860 66946
rect 27804 66052 27860 66894
rect 27916 66948 27972 67006
rect 27916 66882 27972 66892
rect 28028 66724 28084 67452
rect 27804 65986 27860 65996
rect 27916 66668 28084 66724
rect 28252 67172 28308 67182
rect 27916 65602 27972 66668
rect 28252 66274 28308 67116
rect 28364 66388 28420 67900
rect 28364 66322 28420 66332
rect 28252 66222 28254 66274
rect 28306 66222 28308 66274
rect 28252 66210 28308 66222
rect 28140 66162 28196 66174
rect 28140 66110 28142 66162
rect 28194 66110 28196 66162
rect 27916 65550 27918 65602
rect 27970 65550 27972 65602
rect 27916 65538 27972 65550
rect 28028 65716 28084 65726
rect 27692 65438 27694 65490
rect 27746 65438 27748 65490
rect 26908 65212 27188 65268
rect 26908 65044 26964 65054
rect 26908 64594 26964 64988
rect 27020 64932 27076 64942
rect 27020 64838 27076 64876
rect 26908 64542 26910 64594
rect 26962 64542 26964 64594
rect 26908 64530 26964 64542
rect 26796 64094 26798 64146
rect 26850 64094 26852 64146
rect 26796 64082 26852 64094
rect 27132 64148 27188 65212
rect 27468 65044 27524 65054
rect 27468 64818 27524 64988
rect 27468 64766 27470 64818
rect 27522 64766 27524 64818
rect 27468 64754 27524 64766
rect 27132 64082 27188 64092
rect 26516 63868 26628 63924
rect 26460 63858 26516 63868
rect 25900 63250 25956 63756
rect 25900 63198 25902 63250
rect 25954 63198 25956 63250
rect 25900 62692 25956 63198
rect 26348 62914 26404 62926
rect 26348 62862 26350 62914
rect 26402 62862 26404 62914
rect 26348 62692 26404 62862
rect 25956 62636 26180 62692
rect 25900 62626 25956 62636
rect 25564 62578 25732 62580
rect 25564 62526 25566 62578
rect 25618 62526 25732 62578
rect 25564 62524 25732 62526
rect 26124 62578 26180 62636
rect 26348 62626 26404 62636
rect 26124 62526 26126 62578
rect 26178 62526 26180 62578
rect 25564 62514 25620 62524
rect 26124 62514 26180 62526
rect 26572 62580 26628 63868
rect 26684 63922 26740 63934
rect 26684 63870 26686 63922
rect 26738 63870 26740 63922
rect 26684 63812 26740 63870
rect 26908 63924 26964 63934
rect 26908 63830 26964 63868
rect 27132 63924 27188 63934
rect 26684 63746 26740 63756
rect 27132 63252 27188 63868
rect 27356 63924 27412 63934
rect 27692 63924 27748 65438
rect 28028 64708 28084 65660
rect 28140 65492 28196 66110
rect 28140 65426 28196 65436
rect 28364 66162 28420 66174
rect 28364 66110 28366 66162
rect 28418 66110 28420 66162
rect 28364 64932 28420 66110
rect 28364 64866 28420 64876
rect 27804 64706 28084 64708
rect 27804 64654 28030 64706
rect 28082 64654 28084 64706
rect 27804 64652 28084 64654
rect 27804 64146 27860 64652
rect 28028 64642 28084 64652
rect 28252 64820 28308 64830
rect 27804 64094 27806 64146
rect 27858 64094 27860 64146
rect 27804 64082 27860 64094
rect 28252 64036 28308 64764
rect 28252 63970 28308 63980
rect 27356 63922 27748 63924
rect 27356 63870 27358 63922
rect 27410 63870 27748 63922
rect 27356 63868 27748 63870
rect 27356 63858 27412 63868
rect 27244 63252 27300 63262
rect 27132 63250 27300 63252
rect 27132 63198 27246 63250
rect 27298 63198 27300 63250
rect 27132 63196 27300 63198
rect 27244 63186 27300 63196
rect 27692 63250 27748 63868
rect 28476 63364 28532 69244
rect 28812 68964 28868 69358
rect 28812 68898 28868 68908
rect 28700 68516 28756 68526
rect 28700 68422 28756 68460
rect 28812 67956 28868 67966
rect 28812 67862 28868 67900
rect 28588 67172 28644 67182
rect 28588 67078 28644 67116
rect 28812 67060 28868 67070
rect 28700 66948 28756 66958
rect 28588 65716 28644 65726
rect 28588 64146 28644 65660
rect 28588 64094 28590 64146
rect 28642 64094 28644 64146
rect 28588 64082 28644 64094
rect 27692 63198 27694 63250
rect 27746 63198 27748 63250
rect 27580 63140 27636 63150
rect 26796 62916 26852 62926
rect 26796 62822 26852 62860
rect 26684 62580 26740 62590
rect 26572 62578 26740 62580
rect 26572 62526 26686 62578
rect 26738 62526 26740 62578
rect 26572 62524 26740 62526
rect 26684 62514 26740 62524
rect 27580 62578 27636 63084
rect 27692 62916 27748 63198
rect 28364 63308 28532 63364
rect 27692 62850 27748 62860
rect 28252 63140 28308 63150
rect 27580 62526 27582 62578
rect 27634 62526 27636 62578
rect 27580 62514 27636 62526
rect 28252 62578 28308 63084
rect 28252 62526 28254 62578
rect 28306 62526 28308 62578
rect 28252 62514 28308 62526
rect 28364 62580 28420 63308
rect 28700 63252 28756 66892
rect 28812 66498 28868 67004
rect 28924 66724 28980 72156
rect 29148 72604 29316 72660
rect 29148 72100 29204 72604
rect 29596 72548 29652 73892
rect 29708 73330 29764 73342
rect 29708 73278 29710 73330
rect 29762 73278 29764 73330
rect 29708 72884 29764 73278
rect 29820 73330 29876 73342
rect 29820 73278 29822 73330
rect 29874 73278 29876 73330
rect 29820 73220 29876 73278
rect 29820 73154 29876 73164
rect 29708 72818 29764 72828
rect 29036 72044 29204 72100
rect 29260 72492 29652 72548
rect 29820 72660 29876 72670
rect 29036 70196 29092 72044
rect 29148 71764 29204 71774
rect 29148 70420 29204 71708
rect 29260 70532 29316 72492
rect 29596 72322 29652 72334
rect 29596 72270 29598 72322
rect 29650 72270 29652 72322
rect 29372 71874 29428 71886
rect 29372 71822 29374 71874
rect 29426 71822 29428 71874
rect 29372 70980 29428 71822
rect 29372 70914 29428 70924
rect 29484 71652 29540 71662
rect 29372 70532 29428 70542
rect 29260 70476 29372 70532
rect 29372 70466 29428 70476
rect 29148 70364 29316 70420
rect 29148 70196 29204 70206
rect 29036 70194 29204 70196
rect 29036 70142 29150 70194
rect 29202 70142 29204 70194
rect 29036 70140 29204 70142
rect 29036 69412 29092 69422
rect 29036 68626 29092 69356
rect 29036 68574 29038 68626
rect 29090 68574 29092 68626
rect 29036 66948 29092 68574
rect 29148 68628 29204 70140
rect 29148 68180 29204 68572
rect 29148 68114 29204 68124
rect 29260 67396 29316 70364
rect 29484 70418 29540 71596
rect 29596 71540 29652 72270
rect 29596 71474 29652 71484
rect 29708 71428 29764 71438
rect 29596 71204 29652 71214
rect 29596 71110 29652 71148
rect 29708 71202 29764 71372
rect 29708 71150 29710 71202
rect 29762 71150 29764 71202
rect 29708 71092 29764 71150
rect 29708 71026 29764 71036
rect 29820 70868 29876 72604
rect 29484 70366 29486 70418
rect 29538 70366 29540 70418
rect 29484 70354 29540 70366
rect 29708 70812 29876 70868
rect 29932 70978 29988 74172
rect 30044 74564 30100 74574
rect 30044 71762 30100 74508
rect 30268 74564 30324 74574
rect 30268 74116 30324 74508
rect 30268 74022 30324 74060
rect 30268 73108 30324 73118
rect 30156 73106 30324 73108
rect 30156 73054 30270 73106
rect 30322 73054 30324 73106
rect 30156 73052 30324 73054
rect 30156 72548 30212 73052
rect 30268 73042 30324 73052
rect 30268 72884 30324 72894
rect 30268 72770 30324 72828
rect 30268 72718 30270 72770
rect 30322 72718 30324 72770
rect 30268 72706 30324 72718
rect 30156 72492 30324 72548
rect 30268 72212 30324 72492
rect 30380 72322 30436 74844
rect 30492 73948 30548 75740
rect 30604 75348 30660 76526
rect 31724 76578 31780 76636
rect 31724 76526 31726 76578
rect 31778 76526 31780 76578
rect 31724 76514 31780 76526
rect 31836 76580 31892 76860
rect 30940 76356 30996 76366
rect 30940 75682 30996 76300
rect 31276 76242 31332 76254
rect 31276 76190 31278 76242
rect 31330 76190 31332 76242
rect 30940 75630 30942 75682
rect 30994 75630 30996 75682
rect 30940 75618 30996 75630
rect 31052 75794 31108 75806
rect 31052 75742 31054 75794
rect 31106 75742 31108 75794
rect 30604 75282 30660 75292
rect 30828 74900 30884 74910
rect 30828 74806 30884 74844
rect 30604 74340 30660 74350
rect 30604 74226 30660 74284
rect 30604 74174 30606 74226
rect 30658 74174 30660 74226
rect 30604 74162 30660 74174
rect 30940 74002 30996 74014
rect 30940 73950 30942 74002
rect 30994 73950 30996 74002
rect 30492 73892 30660 73948
rect 30492 73556 30548 73566
rect 30492 73442 30548 73500
rect 30492 73390 30494 73442
rect 30546 73390 30548 73442
rect 30492 73108 30548 73390
rect 30492 73042 30548 73052
rect 30604 72996 30660 73892
rect 30940 73332 30996 73950
rect 30940 73266 30996 73276
rect 30380 72270 30382 72322
rect 30434 72270 30436 72322
rect 30380 72258 30436 72270
rect 30492 72660 30548 72670
rect 30268 72146 30324 72156
rect 30044 71710 30046 71762
rect 30098 71710 30100 71762
rect 30044 71698 30100 71710
rect 29932 70926 29934 70978
rect 29986 70926 29988 70978
rect 29596 70308 29652 70318
rect 29596 70214 29652 70252
rect 29372 70194 29428 70206
rect 29372 70142 29374 70194
rect 29426 70142 29428 70194
rect 29372 70084 29428 70142
rect 29708 70084 29764 70812
rect 29820 70308 29876 70318
rect 29820 70214 29876 70252
rect 29372 70028 29764 70084
rect 29372 67956 29428 70028
rect 29932 69412 29988 70926
rect 30044 71540 30100 71550
rect 30044 70084 30100 71484
rect 30156 71316 30212 71326
rect 30156 71202 30212 71260
rect 30156 71150 30158 71202
rect 30210 71150 30212 71202
rect 30156 71138 30212 71150
rect 30380 70980 30436 70990
rect 30380 70756 30436 70924
rect 30380 70690 30436 70700
rect 30492 70308 30548 72604
rect 30604 72324 30660 72940
rect 30940 72772 30996 72782
rect 30604 72258 30660 72268
rect 30716 72546 30772 72558
rect 30716 72494 30718 72546
rect 30770 72494 30772 72546
rect 30604 71764 30660 71774
rect 30716 71764 30772 72494
rect 30828 72546 30884 72558
rect 30828 72494 30830 72546
rect 30882 72494 30884 72546
rect 30828 72436 30884 72494
rect 30828 72370 30884 72380
rect 30660 71708 30772 71764
rect 30604 71670 30660 71708
rect 30492 70242 30548 70252
rect 30044 69860 30100 70028
rect 30044 69794 30100 69804
rect 29820 69356 29988 69412
rect 30156 69524 30212 69534
rect 30156 69410 30212 69468
rect 30156 69358 30158 69410
rect 30210 69358 30212 69410
rect 29708 69186 29764 69198
rect 29708 69134 29710 69186
rect 29762 69134 29764 69186
rect 29708 68852 29764 69134
rect 29708 68786 29764 68796
rect 29820 68180 29876 69356
rect 30156 69346 30212 69358
rect 30268 69412 30324 69422
rect 30044 69300 30100 69310
rect 29932 69188 29988 69226
rect 30044 69206 30100 69244
rect 29932 69122 29988 69132
rect 30044 69076 30100 69086
rect 29932 68964 29988 68974
rect 29932 68402 29988 68908
rect 30044 68738 30100 69020
rect 30044 68686 30046 68738
rect 30098 68686 30100 68738
rect 30044 68674 30100 68686
rect 29932 68350 29934 68402
rect 29986 68350 29988 68402
rect 29932 68338 29988 68350
rect 29820 68124 30100 68180
rect 29596 68068 29652 68078
rect 29596 67974 29652 68012
rect 29372 67890 29428 67900
rect 29820 67956 29876 67966
rect 29708 67618 29764 67630
rect 29708 67566 29710 67618
rect 29762 67566 29764 67618
rect 29260 67340 29540 67396
rect 29148 67172 29204 67182
rect 29260 67172 29316 67340
rect 29204 67116 29316 67172
rect 29372 67172 29428 67182
rect 29148 67106 29204 67116
rect 29260 66948 29316 66958
rect 29036 66946 29316 66948
rect 29036 66894 29262 66946
rect 29314 66894 29316 66946
rect 29036 66892 29316 66894
rect 29260 66882 29316 66892
rect 28924 66658 28980 66668
rect 28812 66446 28814 66498
rect 28866 66446 28868 66498
rect 28812 66434 28868 66446
rect 29372 65828 29428 67116
rect 29484 66612 29540 67340
rect 29596 67060 29652 67070
rect 29596 66966 29652 67004
rect 29708 66948 29764 67566
rect 29708 66882 29764 66892
rect 29484 66556 29764 66612
rect 29596 66386 29652 66398
rect 29596 66334 29598 66386
rect 29650 66334 29652 66386
rect 29596 66276 29652 66334
rect 29596 66210 29652 66220
rect 29372 65762 29428 65772
rect 29708 66162 29764 66556
rect 29820 66500 29876 67900
rect 29932 67732 29988 67742
rect 29932 67638 29988 67676
rect 29932 66500 29988 66510
rect 29820 66498 29988 66500
rect 29820 66446 29934 66498
rect 29986 66446 29988 66498
rect 29820 66444 29988 66446
rect 29708 66110 29710 66162
rect 29762 66110 29764 66162
rect 29708 65716 29764 66110
rect 29484 65490 29540 65502
rect 29484 65438 29486 65490
rect 29538 65438 29540 65490
rect 28812 65378 28868 65390
rect 28812 65326 28814 65378
rect 28866 65326 28868 65378
rect 28812 65156 28868 65326
rect 28812 65090 28868 65100
rect 28924 65380 28980 65390
rect 28924 64148 28980 65324
rect 29484 65380 29540 65438
rect 29708 65490 29764 65660
rect 29708 65438 29710 65490
rect 29762 65438 29764 65490
rect 29708 65426 29764 65438
rect 29932 65828 29988 66444
rect 29484 65314 29540 65324
rect 29820 64820 29876 64830
rect 29932 64820 29988 65772
rect 29876 64764 29988 64820
rect 29820 64688 29876 64764
rect 28924 64016 28980 64092
rect 28812 63252 28868 63262
rect 28700 63250 28868 63252
rect 28700 63198 28814 63250
rect 28866 63198 28868 63250
rect 28700 63196 28868 63198
rect 28812 63140 28868 63196
rect 28812 63074 28868 63084
rect 29932 63140 29988 63150
rect 29932 63046 29988 63084
rect 28364 62466 28420 62524
rect 28364 62414 28366 62466
rect 28418 62414 28420 62466
rect 28364 62402 28420 62414
rect 28476 63028 28532 63038
rect 28028 62354 28084 62366
rect 28028 62302 28030 62354
rect 28082 62302 28084 62354
rect 25340 62244 25396 62254
rect 24892 61954 24948 61964
rect 25116 62020 25172 62030
rect 24556 61618 24612 61628
rect 25004 61908 25060 61918
rect 25004 61682 25060 61852
rect 25004 61630 25006 61682
rect 25058 61630 25060 61682
rect 25004 61618 25060 61630
rect 24108 60958 24110 61010
rect 24162 60958 24164 61010
rect 24108 60946 24164 60958
rect 23660 60114 23828 60116
rect 23660 60062 23662 60114
rect 23714 60062 23828 60114
rect 23660 60060 23828 60062
rect 23660 60050 23716 60060
rect 21308 59378 21364 59388
rect 19516 58930 19572 58940
rect 19628 58884 19684 58894
rect 19516 58660 19572 58670
rect 19404 58658 19572 58660
rect 19404 58606 19518 58658
rect 19570 58606 19572 58658
rect 19404 58604 19572 58606
rect 19516 58594 19572 58604
rect 19628 58548 19684 58828
rect 20076 58548 20132 58558
rect 19628 58546 20132 58548
rect 19628 58494 19630 58546
rect 19682 58494 20078 58546
rect 20130 58494 20132 58546
rect 19628 58492 20132 58494
rect 19628 58482 19684 58492
rect 20076 58482 20132 58492
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19180 57922 19236 57932
rect 18620 56578 18676 56588
rect 19516 57204 19572 57214
rect 17500 50372 18004 50428
rect 16940 36596 16996 36606
rect 17500 36596 17556 50372
rect 19516 48580 19572 57148
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 21868 55412 21924 55422
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 21868 50036 21924 55356
rect 25116 55188 25172 61964
rect 25340 61682 25396 62188
rect 25340 61630 25342 61682
rect 25394 61630 25396 61682
rect 25340 61618 25396 61630
rect 25900 61684 25956 61694
rect 25900 61590 25956 61628
rect 28028 61460 28084 62302
rect 28028 61394 28084 61404
rect 28476 57092 28532 62972
rect 29596 63028 29652 63038
rect 29596 62934 29652 62972
rect 29708 62914 29764 62926
rect 29708 62862 29710 62914
rect 29762 62862 29764 62914
rect 28812 62580 28868 62590
rect 28812 62486 28868 62524
rect 29708 61796 29764 62862
rect 29708 61730 29764 61740
rect 29820 61460 29876 61470
rect 29820 61012 29876 61404
rect 30044 61236 30100 68124
rect 30268 67058 30324 69356
rect 30828 69300 30884 69310
rect 30828 69206 30884 69244
rect 30716 69186 30772 69198
rect 30716 69134 30718 69186
rect 30770 69134 30772 69186
rect 30716 68964 30772 69134
rect 30716 68898 30772 68908
rect 30716 68628 30772 68638
rect 30604 67956 30660 67966
rect 30604 67730 30660 67900
rect 30716 67842 30772 68572
rect 30940 68402 30996 72716
rect 31052 70980 31108 75742
rect 31276 75796 31332 76190
rect 31836 75908 31892 76524
rect 32060 76804 32116 76814
rect 32060 76466 32116 76748
rect 33404 76580 33460 79200
rect 36764 76804 36820 76814
rect 33404 76514 33460 76524
rect 34636 76580 34692 76590
rect 34636 76486 34692 76524
rect 35980 76580 36036 76590
rect 35980 76486 36036 76524
rect 32060 76414 32062 76466
rect 32114 76414 32116 76466
rect 32060 76402 32116 76414
rect 35532 76468 35588 76478
rect 33180 76354 33236 76366
rect 33628 76356 33684 76366
rect 33180 76302 33182 76354
rect 33234 76302 33236 76354
rect 32396 76244 32452 76254
rect 31836 75852 32116 75908
rect 31276 75730 31332 75740
rect 31388 75684 31444 75694
rect 31388 75570 31444 75628
rect 31948 75684 32004 75694
rect 31948 75590 32004 75628
rect 31388 75518 31390 75570
rect 31442 75518 31444 75570
rect 31388 75506 31444 75518
rect 31836 75010 31892 75022
rect 31836 74958 31838 75010
rect 31890 74958 31892 75010
rect 31164 74898 31220 74910
rect 31164 74846 31166 74898
rect 31218 74846 31220 74898
rect 31164 74452 31220 74846
rect 31164 74386 31220 74396
rect 31612 74788 31668 74798
rect 31388 74228 31444 74238
rect 31388 74134 31444 74172
rect 31500 73332 31556 73342
rect 31500 73238 31556 73276
rect 31164 72996 31220 73006
rect 31164 72660 31220 72940
rect 31164 72594 31220 72604
rect 31500 72322 31556 72334
rect 31500 72270 31502 72322
rect 31554 72270 31556 72322
rect 31388 71764 31444 71774
rect 31052 70914 31108 70924
rect 31276 71762 31444 71764
rect 31276 71710 31390 71762
rect 31442 71710 31444 71762
rect 31276 71708 31444 71710
rect 31052 70308 31108 70318
rect 31052 70194 31108 70252
rect 31052 70142 31054 70194
rect 31106 70142 31108 70194
rect 31052 69524 31108 70142
rect 31164 70082 31220 70094
rect 31164 70030 31166 70082
rect 31218 70030 31220 70082
rect 31164 69860 31220 70030
rect 31276 70084 31332 71708
rect 31388 71698 31444 71708
rect 31500 71204 31556 72270
rect 31612 71428 31668 74732
rect 31724 73218 31780 73230
rect 31724 73166 31726 73218
rect 31778 73166 31780 73218
rect 31724 71988 31780 73166
rect 31836 72772 31892 74958
rect 31948 74898 32004 74910
rect 31948 74846 31950 74898
rect 32002 74846 32004 74898
rect 31948 74564 32004 74846
rect 31948 74498 32004 74508
rect 32060 73948 32116 75852
rect 32396 75682 32452 76188
rect 32396 75630 32398 75682
rect 32450 75630 32452 75682
rect 32396 74900 32452 75630
rect 32844 75682 32900 75694
rect 32844 75630 32846 75682
rect 32898 75630 32900 75682
rect 32844 75012 32900 75630
rect 32956 75572 33012 75582
rect 32956 75478 33012 75516
rect 33068 75012 33124 75022
rect 32844 74956 33012 75012
rect 32284 74898 32452 74900
rect 32284 74846 32398 74898
rect 32450 74846 32452 74898
rect 32284 74844 32452 74846
rect 32172 74788 32228 74798
rect 32172 74226 32228 74732
rect 32172 74174 32174 74226
rect 32226 74174 32228 74226
rect 32172 74162 32228 74174
rect 32284 74228 32340 74844
rect 32396 74834 32452 74844
rect 32844 74788 32900 74798
rect 32620 74786 32900 74788
rect 32620 74734 32846 74786
rect 32898 74734 32900 74786
rect 32620 74732 32900 74734
rect 32620 74676 32676 74732
rect 32844 74722 32900 74732
rect 32284 74162 32340 74172
rect 32396 74620 32676 74676
rect 32060 73892 32228 73948
rect 31836 72706 31892 72716
rect 32060 72660 32116 72670
rect 32060 72566 32116 72604
rect 31836 72546 31892 72558
rect 31836 72494 31838 72546
rect 31890 72494 31892 72546
rect 31836 72324 31892 72494
rect 31836 72258 31892 72268
rect 31724 71922 31780 71932
rect 31612 71372 31892 71428
rect 31836 71316 31892 71372
rect 31836 71260 32116 71316
rect 31276 70018 31332 70028
rect 31388 71148 31556 71204
rect 31164 69794 31220 69804
rect 31052 69458 31108 69468
rect 31388 68740 31444 71148
rect 32060 71090 32116 71260
rect 32060 71038 32062 71090
rect 32114 71038 32116 71090
rect 32060 71026 32116 71038
rect 31388 68674 31444 68684
rect 31500 70978 31556 70990
rect 31500 70926 31502 70978
rect 31554 70926 31556 70978
rect 31500 70082 31556 70926
rect 31836 70978 31892 70990
rect 31836 70926 31838 70978
rect 31890 70926 31892 70978
rect 31500 70030 31502 70082
rect 31554 70030 31556 70082
rect 31500 68628 31556 70030
rect 31724 70756 31780 70766
rect 31724 69634 31780 70700
rect 31724 69582 31726 69634
rect 31778 69582 31780 69634
rect 31724 69412 31780 69582
rect 31836 69636 31892 70926
rect 32172 70588 32228 73892
rect 32396 73442 32452 74620
rect 32732 74340 32788 74350
rect 32956 74340 33012 74956
rect 32788 74284 33012 74340
rect 32508 74116 32564 74154
rect 32508 74050 32564 74060
rect 32396 73390 32398 73442
rect 32450 73390 32452 73442
rect 32396 73378 32452 73390
rect 32732 73220 32788 74284
rect 32956 74114 33012 74126
rect 32956 74062 32958 74114
rect 33010 74062 33012 74114
rect 32956 73948 33012 74062
rect 31836 69570 31892 69580
rect 31948 70532 32228 70588
rect 32284 73108 32340 73118
rect 32284 71762 32340 73052
rect 32620 72772 32676 72782
rect 32620 72546 32676 72716
rect 32620 72494 32622 72546
rect 32674 72494 32676 72546
rect 32620 72482 32676 72494
rect 32396 71988 32452 71998
rect 32396 71894 32452 71932
rect 32284 71710 32286 71762
rect 32338 71710 32340 71762
rect 32284 70588 32340 71710
rect 32620 71764 32676 71774
rect 32732 71764 32788 73164
rect 32844 73892 33012 73948
rect 32844 73218 32900 73892
rect 33068 73780 33124 74956
rect 33180 74900 33236 76302
rect 33516 76354 33684 76356
rect 33516 76302 33630 76354
rect 33682 76302 33684 76354
rect 33516 76300 33684 76302
rect 33180 74834 33236 74844
rect 33404 75570 33460 75582
rect 33404 75518 33406 75570
rect 33458 75518 33460 75570
rect 33404 74452 33460 75518
rect 33404 74386 33460 74396
rect 33516 73948 33572 76300
rect 33628 76290 33684 76300
rect 34636 76356 34692 76366
rect 33740 76020 33796 76030
rect 33740 75796 33796 75964
rect 33740 75010 33796 75740
rect 33740 74958 33742 75010
rect 33794 74958 33796 75010
rect 33740 74946 33796 74958
rect 34188 75684 34244 75694
rect 34188 74900 34244 75628
rect 34300 74900 34356 74910
rect 34188 74898 34356 74900
rect 34188 74846 34302 74898
rect 34354 74846 34356 74898
rect 34188 74844 34356 74846
rect 34300 74834 34356 74844
rect 34524 74900 34580 74910
rect 34524 74806 34580 74844
rect 33852 74676 33908 74686
rect 33852 74582 33908 74620
rect 34076 74674 34132 74686
rect 34076 74622 34078 74674
rect 34130 74622 34132 74674
rect 33628 74452 33684 74462
rect 33628 74114 33684 74396
rect 33628 74062 33630 74114
rect 33682 74062 33684 74114
rect 33628 74050 33684 74062
rect 34076 74116 34132 74622
rect 34076 74050 34132 74060
rect 34412 74116 34468 74126
rect 34412 74022 34468 74060
rect 33180 73892 33236 73902
rect 33180 73798 33236 73836
rect 33404 73892 33572 73948
rect 32844 73166 32846 73218
rect 32898 73166 32900 73218
rect 32844 73108 32900 73166
rect 32844 73042 32900 73052
rect 32956 73724 33124 73780
rect 32956 72434 33012 73724
rect 32956 72382 32958 72434
rect 33010 72382 33012 72434
rect 32956 72370 33012 72382
rect 32620 71762 32788 71764
rect 32620 71710 32622 71762
rect 32674 71710 32788 71762
rect 32620 71708 32788 71710
rect 32620 71698 32676 71708
rect 32732 71428 32788 71708
rect 32508 71372 32788 71428
rect 32844 71762 32900 71774
rect 32844 71710 32846 71762
rect 32898 71710 32900 71762
rect 32284 70532 32452 70588
rect 31724 69346 31780 69356
rect 31836 69186 31892 69198
rect 31836 69134 31838 69186
rect 31890 69134 31892 69186
rect 31836 69076 31892 69134
rect 31836 69010 31892 69020
rect 31724 68964 31780 68974
rect 31500 68562 31556 68572
rect 31612 68740 31668 68750
rect 31612 68626 31668 68684
rect 31612 68574 31614 68626
rect 31666 68574 31668 68626
rect 31612 68562 31668 68574
rect 30940 68350 30942 68402
rect 30994 68350 30996 68402
rect 30940 68338 30996 68350
rect 31388 68516 31444 68526
rect 30716 67790 30718 67842
rect 30770 67790 30772 67842
rect 31388 67956 31444 68460
rect 31724 68066 31780 68908
rect 31724 68014 31726 68066
rect 31778 68014 31780 68066
rect 31724 68002 31780 68014
rect 31836 68740 31892 68750
rect 31444 67900 31668 67956
rect 31388 67824 31444 67900
rect 31612 67842 31668 67900
rect 30716 67778 30772 67790
rect 31612 67790 31614 67842
rect 31666 67790 31668 67842
rect 31612 67778 31668 67790
rect 30604 67678 30606 67730
rect 30658 67678 30660 67730
rect 30380 67620 30436 67630
rect 30604 67620 30660 67678
rect 31724 67732 31780 67742
rect 31836 67732 31892 68684
rect 31948 67844 32004 70532
rect 32396 70466 32452 70476
rect 32060 70194 32116 70206
rect 32060 70142 32062 70194
rect 32114 70142 32116 70194
rect 32060 70084 32116 70142
rect 32284 70196 32340 70234
rect 32284 70130 32340 70140
rect 32060 70018 32116 70028
rect 32172 70082 32228 70094
rect 32172 70030 32174 70082
rect 32226 70030 32228 70082
rect 32172 69972 32228 70030
rect 32060 69412 32116 69422
rect 32172 69412 32228 69916
rect 32060 69410 32228 69412
rect 32060 69358 32062 69410
rect 32114 69358 32228 69410
rect 32060 69356 32228 69358
rect 32396 70084 32452 70094
rect 32060 69346 32116 69356
rect 32284 68628 32340 68638
rect 32284 68534 32340 68572
rect 32396 67844 32452 70028
rect 32508 69188 32564 71372
rect 32620 70756 32676 70766
rect 32620 70754 32788 70756
rect 32620 70702 32622 70754
rect 32674 70702 32788 70754
rect 32620 70700 32788 70702
rect 32620 70690 32676 70700
rect 32620 70194 32676 70206
rect 32620 70142 32622 70194
rect 32674 70142 32676 70194
rect 32620 69860 32676 70142
rect 32732 69860 32788 70700
rect 32844 70420 32900 71710
rect 32956 71540 33012 71550
rect 32956 70978 33012 71484
rect 33404 71204 33460 73892
rect 33516 73332 33572 73342
rect 33516 72546 33572 73276
rect 33964 73330 34020 73342
rect 33964 73278 33966 73330
rect 34018 73278 34020 73330
rect 33740 73218 33796 73230
rect 33740 73166 33742 73218
rect 33794 73166 33796 73218
rect 33740 73108 33796 73166
rect 33740 73042 33796 73052
rect 33964 73220 34020 73278
rect 34636 73220 34692 76300
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 34972 75684 35028 75694
rect 33964 72770 34020 73164
rect 33964 72718 33966 72770
rect 34018 72718 34020 72770
rect 33964 72706 34020 72718
rect 34524 73218 34692 73220
rect 34524 73166 34638 73218
rect 34690 73166 34692 73218
rect 34524 73164 34692 73166
rect 33516 72494 33518 72546
rect 33570 72494 33572 72546
rect 33516 72482 33572 72494
rect 33628 72322 33684 72334
rect 33628 72270 33630 72322
rect 33682 72270 33684 72322
rect 33628 71652 33684 72270
rect 33852 72324 33908 72334
rect 34188 72324 34244 72334
rect 34524 72324 34580 73164
rect 34636 73154 34692 73164
rect 34860 75682 35028 75684
rect 34860 75630 34974 75682
rect 35026 75630 35028 75682
rect 34860 75628 35028 75630
rect 34860 74788 34916 75628
rect 34972 75618 35028 75628
rect 35420 75124 35476 75134
rect 35532 75124 35588 76412
rect 35420 75122 35588 75124
rect 35420 75070 35422 75122
rect 35474 75070 35588 75122
rect 35420 75068 35588 75070
rect 35644 76356 35700 76366
rect 36540 76356 36596 76366
rect 35644 76354 35812 76356
rect 35644 76302 35646 76354
rect 35698 76302 35812 76354
rect 35644 76300 35812 76302
rect 35644 75684 35700 76300
rect 35756 76244 35812 76300
rect 35756 76178 35812 76188
rect 36540 75794 36596 76300
rect 36764 76356 36820 76748
rect 37548 76692 37604 76702
rect 37772 76692 37828 79200
rect 38668 77812 38724 77822
rect 37548 76690 37828 76692
rect 37548 76638 37550 76690
rect 37602 76638 37828 76690
rect 37548 76636 37828 76638
rect 37548 76626 37604 76636
rect 37772 76580 37828 76636
rect 37772 76514 37828 76524
rect 37884 77700 37940 77710
rect 37100 76356 37156 76366
rect 36764 76290 36820 76300
rect 36988 76354 37156 76356
rect 36988 76302 37102 76354
rect 37154 76302 37156 76354
rect 36988 76300 37156 76302
rect 36540 75742 36542 75794
rect 36594 75742 36596 75794
rect 36540 75730 36596 75742
rect 35644 75124 35700 75628
rect 36092 75572 36148 75582
rect 36092 75478 36148 75516
rect 35756 75460 35812 75470
rect 35756 75458 36036 75460
rect 35756 75406 35758 75458
rect 35810 75406 36036 75458
rect 35756 75404 36036 75406
rect 35756 75394 35812 75404
rect 35868 75124 35924 75134
rect 35644 75122 35924 75124
rect 35644 75070 35870 75122
rect 35922 75070 35924 75122
rect 35644 75068 35924 75070
rect 35420 74900 35476 75068
rect 35868 75058 35924 75068
rect 35420 74834 35476 74844
rect 34860 74564 34916 74732
rect 34748 72996 34804 73006
rect 34636 72770 34692 72782
rect 34636 72718 34638 72770
rect 34690 72718 34692 72770
rect 34636 72658 34692 72718
rect 34636 72606 34638 72658
rect 34690 72606 34692 72658
rect 34636 72594 34692 72606
rect 33852 72230 33908 72268
rect 33964 72322 34580 72324
rect 33964 72270 34190 72322
rect 34242 72270 34580 72322
rect 33964 72268 34580 72270
rect 34748 72324 34804 72940
rect 33852 71876 33908 71886
rect 33852 71782 33908 71820
rect 33964 71652 34020 72268
rect 34188 72258 34244 72268
rect 34076 71988 34132 71998
rect 34076 71986 34356 71988
rect 34076 71934 34078 71986
rect 34130 71934 34356 71986
rect 34076 71932 34356 71934
rect 34076 71922 34132 71932
rect 33628 71596 34020 71652
rect 33404 71138 33460 71148
rect 32956 70926 32958 70978
rect 33010 70926 33012 70978
rect 32956 70914 33012 70926
rect 33404 70980 33460 70990
rect 33740 70980 33796 70990
rect 33404 70886 33460 70924
rect 33516 70978 33796 70980
rect 33516 70926 33742 70978
rect 33794 70926 33796 70978
rect 33516 70924 33796 70926
rect 32844 70354 32900 70364
rect 33292 70756 33348 70766
rect 32732 69804 32900 69860
rect 32620 69300 32676 69804
rect 32732 69636 32788 69646
rect 32732 69542 32788 69580
rect 32844 69412 32900 69804
rect 32844 69356 33012 69412
rect 32620 69234 32676 69244
rect 32844 69242 32900 69254
rect 32508 68852 32564 69132
rect 32508 68786 32564 68796
rect 32732 69186 32788 69198
rect 32732 69134 32734 69186
rect 32786 69134 32788 69186
rect 32620 68626 32676 68638
rect 32620 68574 32622 68626
rect 32674 68574 32676 68626
rect 32620 68516 32676 68574
rect 32620 68450 32676 68460
rect 31948 67788 32228 67844
rect 31724 67730 31892 67732
rect 31724 67678 31726 67730
rect 31778 67678 31892 67730
rect 31724 67676 31892 67678
rect 30380 67618 30548 67620
rect 30380 67566 30382 67618
rect 30434 67566 30548 67618
rect 30380 67564 30548 67566
rect 30604 67564 30772 67620
rect 30380 67554 30436 67564
rect 30268 67006 30270 67058
rect 30322 67006 30324 67058
rect 30268 66994 30324 67006
rect 30492 67060 30548 67564
rect 30604 67060 30660 67070
rect 30492 67058 30660 67060
rect 30492 67006 30606 67058
rect 30658 67006 30660 67058
rect 30492 67004 30660 67006
rect 30604 66994 30660 67004
rect 30716 66836 30772 67564
rect 31388 67282 31444 67294
rect 31388 67230 31390 67282
rect 31442 67230 31444 67282
rect 31388 67172 31444 67230
rect 31612 67284 31668 67294
rect 31724 67284 31780 67676
rect 31612 67282 31780 67284
rect 31612 67230 31614 67282
rect 31666 67230 31780 67282
rect 31612 67228 31780 67230
rect 31948 67620 32004 67630
rect 31948 67282 32004 67564
rect 31948 67230 31950 67282
rect 32002 67230 32004 67282
rect 31612 67218 31668 67228
rect 31388 67106 31444 67116
rect 31276 67060 31332 67070
rect 31276 66966 31332 67004
rect 30604 66780 30772 66836
rect 30604 66386 30660 66780
rect 30604 66334 30606 66386
rect 30658 66334 30660 66386
rect 30604 66322 30660 66334
rect 31276 66724 31332 66734
rect 31276 66274 31332 66668
rect 31948 66724 32004 67230
rect 31948 66658 32004 66668
rect 32060 66834 32116 66846
rect 32060 66782 32062 66834
rect 32114 66782 32116 66834
rect 31276 66222 31278 66274
rect 31330 66222 31332 66274
rect 30604 65828 30660 65838
rect 30492 65716 30548 65726
rect 30492 65622 30548 65660
rect 30380 65604 30436 65614
rect 30268 65492 30324 65502
rect 30268 65398 30324 65436
rect 30268 64820 30324 64830
rect 30380 64820 30436 65548
rect 30604 65602 30660 65772
rect 31052 65716 31108 65726
rect 31052 65622 31108 65660
rect 30604 65550 30606 65602
rect 30658 65550 30660 65602
rect 30604 65538 30660 65550
rect 31276 65604 31332 66222
rect 31276 65538 31332 65548
rect 31500 66388 31556 66398
rect 32060 66388 32116 66782
rect 31500 66386 32116 66388
rect 31500 66334 31502 66386
rect 31554 66334 32062 66386
rect 32114 66334 32116 66386
rect 31500 66332 32116 66334
rect 31500 65380 31556 66332
rect 32060 66322 32116 66332
rect 31500 65314 31556 65324
rect 30268 64818 30436 64820
rect 30268 64766 30270 64818
rect 30322 64766 30436 64818
rect 30268 64764 30436 64766
rect 30268 64754 30324 64764
rect 30044 61170 30100 61180
rect 30380 62916 30436 62926
rect 30380 61012 30436 62860
rect 30940 61012 30996 61022
rect 29820 61010 30324 61012
rect 29820 60958 29822 61010
rect 29874 60958 30324 61010
rect 29820 60956 30324 60958
rect 29820 60946 29876 60956
rect 30268 60898 30324 60956
rect 30380 61010 30996 61012
rect 30380 60958 30382 61010
rect 30434 60958 30942 61010
rect 30994 60958 30996 61010
rect 30380 60956 30996 60958
rect 30380 60946 30436 60956
rect 30940 60946 30996 60956
rect 30268 60846 30270 60898
rect 30322 60846 30324 60898
rect 30268 60834 30324 60846
rect 30380 60562 30436 60574
rect 30380 60510 30382 60562
rect 30434 60510 30436 60562
rect 30380 60340 30436 60510
rect 30380 60274 30436 60284
rect 28476 57026 28532 57036
rect 28812 56644 28868 56654
rect 25116 54964 25172 55132
rect 27804 56308 27860 56318
rect 25116 54898 25172 54908
rect 26012 54964 26068 54974
rect 21868 49970 21924 49980
rect 23212 50036 23268 50046
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19516 48514 19572 48524
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 16940 36594 17556 36596
rect 16940 36542 16942 36594
rect 16994 36542 17556 36594
rect 16940 36540 17556 36542
rect 16940 36530 16996 36540
rect 17500 36482 17556 36540
rect 17500 36430 17502 36482
rect 17554 36430 17556 36482
rect 17500 6804 17556 36430
rect 17612 36708 17668 36718
rect 17612 36260 17668 36652
rect 17612 36194 17668 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 17500 6738 17556 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 18620 6020 18676 6030
rect 18620 5906 18676 5964
rect 19628 6020 19684 6030
rect 19628 5926 19684 5964
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5842 18676 5854
rect 18172 5796 18228 5806
rect 18172 5702 18228 5740
rect 18844 5796 18900 5806
rect 16716 5282 16772 5292
rect 18844 5682 18900 5740
rect 18844 5630 18846 5682
rect 18898 5630 18900 5682
rect 18844 5124 18900 5630
rect 19180 5684 19236 5694
rect 19180 5682 19572 5684
rect 19180 5630 19182 5682
rect 19234 5630 19572 5682
rect 19180 5628 19572 5630
rect 19180 5618 19236 5628
rect 18844 5058 18900 5068
rect 15148 4340 15204 4350
rect 15036 4338 15204 4340
rect 15036 4286 15150 4338
rect 15202 4286 15204 4338
rect 15036 4284 15204 4286
rect 11564 3502 11566 3554
rect 11618 3502 11620 3554
rect 11564 3490 11620 3502
rect 11676 3668 11732 3678
rect 11676 800 11732 3612
rect 12236 3668 12292 3678
rect 12236 3574 12292 3612
rect 15148 3668 15204 4284
rect 15372 4338 15428 4508
rect 16604 4452 16660 4462
rect 16604 4358 16660 4396
rect 17500 4452 17556 4462
rect 19516 4452 19572 5628
rect 22764 5236 22820 5246
rect 23212 5236 23268 49980
rect 22764 5234 23268 5236
rect 22764 5182 22766 5234
rect 22818 5182 23214 5234
rect 23266 5182 23268 5234
rect 22764 5180 23268 5182
rect 22764 5170 22820 5180
rect 23212 5170 23268 5180
rect 26012 5236 26068 54908
rect 26012 5170 26068 5180
rect 22204 5124 22260 5134
rect 22204 5030 22260 5068
rect 23436 5124 23492 5134
rect 23436 5030 23492 5068
rect 26796 5124 26852 5134
rect 23772 5012 23828 5022
rect 24332 5012 24388 5022
rect 23772 5010 24388 5012
rect 23772 4958 23774 5010
rect 23826 4958 24334 5010
rect 24386 4958 24388 5010
rect 23772 4956 24388 4958
rect 23772 4946 23828 4956
rect 24332 4946 24388 4956
rect 24668 4900 24724 4910
rect 24668 4806 24724 4844
rect 26012 4900 26068 4910
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4452 19684 4462
rect 19516 4450 19684 4452
rect 19516 4398 19630 4450
rect 19682 4398 19684 4450
rect 19516 4396 19684 4398
rect 15372 4286 15374 4338
rect 15426 4286 15428 4338
rect 15372 4274 15428 4286
rect 15708 4340 15764 4350
rect 16268 4340 16324 4350
rect 15708 4338 16324 4340
rect 15708 4286 15710 4338
rect 15762 4286 16270 4338
rect 16322 4286 16324 4338
rect 15708 4284 16324 4286
rect 15708 4274 15764 4284
rect 16268 4274 16324 4284
rect 15148 3602 15204 3612
rect 16044 3668 16100 3678
rect 16044 3574 16100 3612
rect 16380 3668 16436 3678
rect 16380 800 16436 3612
rect 17500 3554 17556 4396
rect 19628 4386 19684 4396
rect 19964 4452 20020 4462
rect 19964 4358 20020 4396
rect 21420 4452 21476 4462
rect 18172 3668 18228 3678
rect 18172 3574 18228 3612
rect 21084 3668 21140 3678
rect 17500 3502 17502 3554
rect 17554 3502 17556 3554
rect 17500 3490 17556 3502
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21084 800 21140 3612
rect 21420 3554 21476 4396
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 25788 3668 25844 3678
rect 21420 3502 21422 3554
rect 21474 3502 21476 3554
rect 21420 3490 21476 3502
rect 25788 800 25844 3612
rect 26012 3554 26068 4844
rect 26796 4562 26852 5068
rect 26796 4510 26798 4562
rect 26850 4510 26852 4562
rect 26796 4498 26852 4510
rect 27244 4564 27300 4574
rect 27804 4564 27860 56252
rect 28812 55524 28868 56588
rect 28812 55298 28868 55468
rect 28812 55246 28814 55298
rect 28866 55246 28868 55298
rect 28812 55234 28868 55246
rect 29596 55524 29652 55534
rect 29596 55298 29652 55468
rect 32172 55468 32228 67788
rect 32396 67842 32676 67844
rect 32396 67790 32398 67842
rect 32450 67790 32676 67842
rect 32396 67788 32676 67790
rect 32396 67778 32452 67788
rect 32508 67620 32564 67630
rect 32508 67526 32564 67564
rect 32620 67620 32676 67788
rect 32732 67842 32788 69134
rect 32844 69190 32846 69242
rect 32898 69190 32900 69242
rect 32844 68964 32900 69190
rect 32956 69076 33012 69356
rect 32956 69020 33236 69076
rect 32844 68898 32900 68908
rect 32956 68852 33012 68862
rect 32956 68758 33012 68796
rect 32844 68740 32900 68750
rect 32844 68646 32900 68684
rect 32732 67790 32734 67842
rect 32786 67790 32788 67842
rect 32732 67778 32788 67790
rect 33068 67620 33124 67630
rect 32620 67618 33124 67620
rect 32620 67566 33070 67618
rect 33122 67566 33124 67618
rect 32620 67564 33124 67566
rect 32396 67172 32452 67182
rect 32396 67078 32452 67116
rect 32620 66834 32676 67564
rect 33068 67554 33124 67564
rect 32844 67172 32900 67182
rect 32844 67078 32900 67116
rect 32620 66782 32622 66834
rect 32674 66782 32676 66834
rect 32620 66770 32676 66782
rect 33180 56868 33236 69020
rect 33292 62020 33348 70700
rect 33516 70194 33572 70924
rect 33740 70914 33796 70924
rect 33628 70756 33684 70766
rect 33628 70754 33908 70756
rect 33628 70702 33630 70754
rect 33682 70702 33908 70754
rect 33628 70700 33908 70702
rect 33628 70690 33684 70700
rect 33740 70420 33796 70430
rect 33740 70326 33796 70364
rect 33516 70142 33518 70194
rect 33570 70142 33572 70194
rect 33516 69972 33572 70142
rect 33516 69906 33572 69916
rect 33852 70194 33908 70700
rect 33852 70142 33854 70194
rect 33906 70142 33908 70194
rect 33516 69636 33572 69646
rect 33516 69542 33572 69580
rect 33404 69412 33460 69422
rect 33404 69318 33460 69356
rect 33516 69300 33572 69310
rect 33516 68740 33572 69244
rect 33852 68852 33908 70142
rect 33964 69412 34020 71596
rect 34188 71762 34244 71774
rect 34188 71710 34190 71762
rect 34242 71710 34244 71762
rect 34188 70754 34244 71710
rect 34188 70702 34190 70754
rect 34242 70702 34244 70754
rect 34076 70194 34132 70206
rect 34076 70142 34078 70194
rect 34130 70142 34132 70194
rect 34076 69636 34132 70142
rect 34076 69570 34132 69580
rect 34076 69412 34132 69422
rect 33964 69356 34076 69412
rect 34076 69318 34132 69356
rect 33852 68786 33908 68796
rect 33964 69188 34020 69198
rect 33964 68850 34020 69132
rect 33964 68798 33966 68850
rect 34018 68798 34020 68850
rect 33964 68786 34020 68798
rect 33516 68646 33572 68684
rect 34188 68180 34244 70702
rect 34188 68114 34244 68124
rect 34300 71652 34356 71932
rect 34636 71652 34692 71662
rect 34300 71650 34692 71652
rect 34300 71598 34638 71650
rect 34690 71598 34692 71650
rect 34300 71596 34692 71598
rect 33964 67732 34020 67742
rect 33964 67638 34020 67676
rect 33516 67618 33572 67630
rect 33516 67566 33518 67618
rect 33570 67566 33572 67618
rect 33516 66948 33572 67566
rect 33516 66882 33572 66892
rect 34300 63252 34356 71596
rect 34636 71586 34692 71596
rect 34636 70980 34692 70990
rect 34636 70886 34692 70924
rect 34636 70084 34692 70094
rect 34636 69990 34692 70028
rect 34524 69524 34580 69534
rect 34748 69524 34804 72268
rect 34524 69522 34804 69524
rect 34524 69470 34526 69522
rect 34578 69470 34804 69522
rect 34524 69468 34804 69470
rect 34860 70420 34916 74508
rect 34972 74786 35028 74798
rect 34972 74734 34974 74786
rect 35026 74734 35028 74786
rect 34972 74116 35028 74734
rect 35980 74676 36036 75404
rect 36988 75124 37044 76300
rect 37100 76290 37156 76300
rect 37548 76132 37604 76142
rect 37324 75908 37380 75918
rect 36316 74786 36372 74798
rect 36316 74734 36318 74786
rect 36370 74734 36372 74786
rect 36316 74676 36372 74734
rect 36764 74788 36820 74798
rect 36764 74694 36820 74732
rect 35980 74620 36260 74676
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 36092 74452 36148 74462
rect 34972 74050 35028 74060
rect 35196 74228 35252 74238
rect 35196 74114 35252 74172
rect 35196 74062 35198 74114
rect 35250 74062 35252 74114
rect 35196 73948 35252 74062
rect 35980 74116 36036 74126
rect 35980 74022 36036 74060
rect 34972 73892 35252 73948
rect 34972 72770 35028 73892
rect 35196 73556 35252 73892
rect 35644 73780 35700 73790
rect 35532 73556 35588 73566
rect 35196 73554 35588 73556
rect 35196 73502 35534 73554
rect 35586 73502 35588 73554
rect 35196 73500 35588 73502
rect 35084 73218 35140 73230
rect 35084 73166 35086 73218
rect 35138 73166 35140 73218
rect 35084 73108 35140 73166
rect 35084 73042 35140 73052
rect 35532 73106 35588 73500
rect 35532 73054 35534 73106
rect 35586 73054 35588 73106
rect 35532 73042 35588 73054
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 34972 72718 34974 72770
rect 35026 72718 35028 72770
rect 34972 72706 35028 72718
rect 35644 72772 35700 73724
rect 35980 73218 36036 73230
rect 35980 73166 35982 73218
rect 36034 73166 36036 73218
rect 35980 73106 36036 73166
rect 35980 73054 35982 73106
rect 36034 73054 36036 73106
rect 35980 73042 36036 73054
rect 35644 72658 35700 72716
rect 35644 72606 35646 72658
rect 35698 72606 35700 72658
rect 35644 72594 35700 72606
rect 35980 72884 36036 72894
rect 35980 72436 36036 72828
rect 35980 72342 36036 72380
rect 35084 72324 35140 72334
rect 35084 72230 35140 72268
rect 35084 71876 35140 71886
rect 35084 71782 35140 71820
rect 35532 71876 35588 71886
rect 35532 71782 35588 71820
rect 35980 71650 36036 71662
rect 35980 71598 35982 71650
rect 36034 71598 36036 71650
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 71204 35252 71214
rect 35196 71090 35252 71148
rect 35980 71204 36036 71598
rect 35980 71138 36036 71148
rect 35196 71038 35198 71090
rect 35250 71038 35252 71090
rect 35196 71026 35252 71038
rect 35532 71092 35588 71102
rect 35532 70998 35588 71036
rect 35980 70756 36036 70766
rect 34860 69522 34916 70364
rect 35532 70754 36036 70756
rect 35532 70702 35982 70754
rect 36034 70702 36036 70754
rect 35532 70700 36036 70702
rect 35084 70308 35140 70318
rect 35084 70214 35140 70252
rect 35532 70084 35588 70700
rect 35980 70690 36036 70700
rect 35644 70420 35700 70430
rect 36092 70420 36148 74396
rect 35644 70418 36148 70420
rect 35644 70366 35646 70418
rect 35698 70366 36148 70418
rect 35644 70364 36148 70366
rect 35644 70354 35700 70364
rect 35532 70018 35588 70028
rect 35756 70196 35812 70206
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 34860 69470 34862 69522
rect 34914 69470 34916 69522
rect 34524 69458 34580 69468
rect 34860 69458 34916 69470
rect 35308 69636 35364 69646
rect 35308 69522 35364 69580
rect 35308 69470 35310 69522
rect 35362 69470 35364 69522
rect 35308 69458 35364 69470
rect 35756 69522 35812 70140
rect 35756 69470 35758 69522
rect 35810 69470 35812 69522
rect 35756 69458 35812 69470
rect 35980 70082 36036 70094
rect 35980 70030 35982 70082
rect 36034 70030 36036 70082
rect 35980 69970 36036 70030
rect 35980 69918 35982 69970
rect 36034 69918 36036 69970
rect 35532 68852 35588 68862
rect 34524 68740 34580 68750
rect 34412 68516 34468 68526
rect 34412 67844 34468 68460
rect 34412 67778 34468 67788
rect 34412 67620 34468 67630
rect 34524 67620 34580 68684
rect 34860 68514 34916 68526
rect 34860 68462 34862 68514
rect 34914 68462 34916 68514
rect 34860 68180 34916 68462
rect 35308 68514 35364 68526
rect 35308 68462 35310 68514
rect 35362 68462 35364 68514
rect 35308 68404 35364 68462
rect 35308 68338 35364 68348
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 34860 68114 34916 68124
rect 34468 67564 34580 67620
rect 34412 67488 34468 67564
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35532 66500 35588 68796
rect 35980 67508 36036 69918
rect 36204 69412 36260 74620
rect 36316 74610 36372 74620
rect 36540 74340 36596 74350
rect 36540 74228 36596 74284
rect 36764 74228 36820 74238
rect 36988 74228 37044 75068
rect 36540 74226 37044 74228
rect 36540 74174 36766 74226
rect 36818 74174 37044 74226
rect 36540 74172 37044 74174
rect 37100 75906 37380 75908
rect 37100 75854 37326 75906
rect 37378 75854 37380 75906
rect 37100 75852 37380 75854
rect 36316 73890 36372 73902
rect 36316 73838 36318 73890
rect 36370 73838 36372 73890
rect 36316 73108 36372 73838
rect 36428 73780 36484 73790
rect 36428 73554 36484 73724
rect 36428 73502 36430 73554
rect 36482 73502 36484 73554
rect 36428 73490 36484 73502
rect 36316 73042 36372 73052
rect 36428 72660 36484 72670
rect 36428 72212 36484 72604
rect 36428 72146 36484 72156
rect 35980 67442 36036 67452
rect 36092 69356 36260 69412
rect 36316 72100 36372 72110
rect 35532 66434 35588 66444
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 34300 63186 34356 63196
rect 33292 61954 33348 61964
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 33180 56802 33236 56812
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 32172 55412 32676 55468
rect 29596 55246 29598 55298
rect 29650 55246 29652 55298
rect 29596 55234 29652 55246
rect 29932 55076 29988 55086
rect 29932 54982 29988 55020
rect 32620 41972 32676 55412
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 36092 52052 36148 69356
rect 36204 69188 36260 69198
rect 36316 69188 36372 72044
rect 36428 71650 36484 71662
rect 36428 71598 36430 71650
rect 36482 71598 36484 71650
rect 36428 71538 36484 71598
rect 36428 71486 36430 71538
rect 36482 71486 36484 71538
rect 36428 71474 36484 71486
rect 36428 71092 36484 71102
rect 36540 71092 36596 74172
rect 36764 74162 36820 74172
rect 36876 73444 36932 73454
rect 36876 73350 36932 73388
rect 36876 71988 36932 71998
rect 36876 71652 36932 71932
rect 36876 71586 36932 71596
rect 36428 71090 36596 71092
rect 36428 71038 36430 71090
rect 36482 71038 36596 71090
rect 36428 71036 36596 71038
rect 36652 71538 36708 71550
rect 36652 71486 36654 71538
rect 36706 71486 36708 71538
rect 36428 71026 36484 71036
rect 36428 70420 36484 70430
rect 36428 70326 36484 70364
rect 36652 69970 36708 71486
rect 37100 70980 37156 75852
rect 37324 75842 37380 75852
rect 37436 75458 37492 75470
rect 37436 75406 37438 75458
rect 37490 75406 37492 75458
rect 37212 74788 37268 74798
rect 37212 74694 37268 74732
rect 37324 74338 37380 74350
rect 37324 74286 37326 74338
rect 37378 74286 37380 74338
rect 37324 73948 37380 74286
rect 37436 74228 37492 75406
rect 37436 74162 37492 74172
rect 37548 75460 37604 76076
rect 37884 75684 37940 77644
rect 38332 76916 38388 76926
rect 37996 76354 38052 76366
rect 37996 76302 37998 76354
rect 38050 76302 38052 76354
rect 37996 75906 38052 76302
rect 37996 75854 37998 75906
rect 38050 75854 38052 75906
rect 37996 75842 38052 75854
rect 38220 75908 38276 75918
rect 37884 75628 38052 75684
rect 37884 75460 37940 75470
rect 37548 75458 37940 75460
rect 37548 75406 37886 75458
rect 37938 75406 37940 75458
rect 37548 75404 37940 75406
rect 37548 74674 37604 75404
rect 37884 75394 37940 75404
rect 37660 74788 37716 74798
rect 37660 74694 37716 74732
rect 37548 74622 37550 74674
rect 37602 74622 37604 74674
rect 37100 70914 37156 70924
rect 37212 73892 37380 73948
rect 37436 74002 37492 74014
rect 37436 73950 37438 74002
rect 37490 73950 37492 74002
rect 37436 73948 37492 73950
rect 37548 73948 37604 74622
rect 37884 74228 37940 74238
rect 37884 74134 37940 74172
rect 37436 73892 37604 73948
rect 37212 71092 37268 73892
rect 37324 73556 37380 73566
rect 37324 73462 37380 73500
rect 37436 72772 37492 73892
rect 37324 72716 37492 72772
rect 37772 73218 37828 73230
rect 37772 73166 37774 73218
rect 37826 73166 37828 73218
rect 37324 71986 37380 72716
rect 37324 71934 37326 71986
rect 37378 71934 37380 71986
rect 37324 71922 37380 71934
rect 37436 72322 37492 72334
rect 37436 72270 37438 72322
rect 37490 72270 37492 72322
rect 37436 71538 37492 72270
rect 37772 72100 37828 73166
rect 37884 72660 37940 72670
rect 37996 72660 38052 75628
rect 38220 75236 38276 75852
rect 38332 75794 38388 76860
rect 38332 75742 38334 75794
rect 38386 75742 38388 75794
rect 38332 75730 38388 75742
rect 38220 75180 38388 75236
rect 38108 74786 38164 74798
rect 38108 74734 38110 74786
rect 38162 74734 38164 74786
rect 38108 74338 38164 74734
rect 38108 74286 38110 74338
rect 38162 74286 38164 74338
rect 38108 74274 38164 74286
rect 38332 74226 38388 75180
rect 38556 75124 38612 75134
rect 38556 75030 38612 75068
rect 38668 74676 38724 77756
rect 40124 77588 40180 77598
rect 39900 76692 39956 76702
rect 39900 76598 39956 76636
rect 39004 76580 39060 76590
rect 39004 76486 39060 76524
rect 38780 76356 38836 76366
rect 38780 75794 38836 76300
rect 38780 75742 38782 75794
rect 38834 75742 38836 75794
rect 38780 75730 38836 75742
rect 40124 75794 40180 77532
rect 40908 77476 40964 77486
rect 40908 76690 40964 77420
rect 40908 76638 40910 76690
rect 40962 76638 40964 76690
rect 40908 76626 40964 76638
rect 41916 76692 41972 76702
rect 42140 76692 42196 79200
rect 41916 76690 42196 76692
rect 41916 76638 41918 76690
rect 41970 76638 42196 76690
rect 41916 76636 42196 76638
rect 41916 76626 41972 76636
rect 42140 76580 42196 76636
rect 42140 76514 42196 76524
rect 43372 76580 43428 76590
rect 43372 76486 43428 76524
rect 46508 76580 46564 79200
rect 48860 78036 48916 78046
rect 46508 76514 46564 76524
rect 47628 76580 47684 76590
rect 47628 76486 47684 76524
rect 48748 76580 48804 76590
rect 48748 76486 48804 76524
rect 40124 75742 40126 75794
rect 40178 75742 40180 75794
rect 40124 75730 40180 75742
rect 41356 76354 41412 76366
rect 41356 76302 41358 76354
rect 41410 76302 41412 76354
rect 39452 75684 39508 75694
rect 39228 75458 39284 75470
rect 39228 75406 39230 75458
rect 39282 75406 39284 75458
rect 39228 75348 39284 75406
rect 39228 75282 39284 75292
rect 39452 75122 39508 75628
rect 39452 75070 39454 75122
rect 39506 75070 39508 75122
rect 39452 75058 39508 75070
rect 39676 75458 39732 75470
rect 39676 75406 39678 75458
rect 39730 75406 39732 75458
rect 39004 74786 39060 74798
rect 39004 74734 39006 74786
rect 39058 74734 39060 74786
rect 38668 74620 38836 74676
rect 38332 74174 38334 74226
rect 38386 74174 38388 74226
rect 38332 74162 38388 74174
rect 38668 74338 38724 74350
rect 38668 74286 38670 74338
rect 38722 74286 38724 74338
rect 38668 73892 38724 74286
rect 38780 74226 38836 74620
rect 39004 74674 39060 74734
rect 39004 74622 39006 74674
rect 39058 74622 39060 74674
rect 39004 74610 39060 74622
rect 38780 74174 38782 74226
rect 38834 74174 38836 74226
rect 38780 74162 38836 74174
rect 38668 73826 38724 73836
rect 39228 73890 39284 73902
rect 39676 73892 39732 75406
rect 40572 75460 40628 75470
rect 41020 75460 41076 75470
rect 41356 75460 41412 76302
rect 42364 76354 42420 76366
rect 42364 76302 42366 76354
rect 42418 76302 42420 76354
rect 40572 75458 41412 75460
rect 40572 75406 40574 75458
rect 40626 75406 41022 75458
rect 41074 75406 41412 75458
rect 40572 75404 41412 75406
rect 41468 75458 41524 75470
rect 41468 75406 41470 75458
rect 41522 75406 41524 75458
rect 39900 74786 39956 74798
rect 40348 74788 40404 74798
rect 40572 74788 40628 75404
rect 41020 75394 41076 75404
rect 41468 75012 41524 75406
rect 41356 74956 41524 75012
rect 41916 75458 41972 75470
rect 41916 75406 41918 75458
rect 41970 75406 41972 75458
rect 39900 74734 39902 74786
rect 39954 74734 39956 74786
rect 39900 74338 39956 74734
rect 39900 74286 39902 74338
rect 39954 74286 39956 74338
rect 39900 74274 39956 74286
rect 40124 74786 40628 74788
rect 40124 74734 40350 74786
rect 40402 74734 40628 74786
rect 40124 74732 40628 74734
rect 40796 74786 40852 74798
rect 40796 74734 40798 74786
rect 40850 74734 40852 74786
rect 40124 73892 40180 74732
rect 40348 74722 40404 74732
rect 39228 73838 39230 73890
rect 39282 73838 39284 73890
rect 38220 73220 38276 73230
rect 37884 72658 38052 72660
rect 37884 72606 37886 72658
rect 37938 72606 38052 72658
rect 37884 72604 38052 72606
rect 38108 73218 38276 73220
rect 38108 73166 38222 73218
rect 38274 73166 38276 73218
rect 38108 73164 38276 73166
rect 37884 72594 37940 72604
rect 37772 72034 37828 72044
rect 37436 71486 37438 71538
rect 37490 71486 37492 71538
rect 37436 71474 37492 71486
rect 37772 71764 37828 71774
rect 37436 71092 37492 71102
rect 37212 71090 37492 71092
rect 37212 71038 37438 71090
rect 37490 71038 37492 71090
rect 37212 71036 37492 71038
rect 37212 70532 37268 71036
rect 37436 71026 37492 71036
rect 37772 70644 37828 71708
rect 37772 70578 37828 70588
rect 37884 70754 37940 70766
rect 37884 70702 37886 70754
rect 37938 70702 37940 70754
rect 37212 70466 37268 70476
rect 36988 70196 37044 70206
rect 36988 70102 37044 70140
rect 37324 70196 37380 70206
rect 37324 70102 37380 70140
rect 36652 69918 36654 69970
rect 36706 69918 36708 69970
rect 36652 69906 36708 69918
rect 36204 69186 36372 69188
rect 36204 69134 36206 69186
rect 36258 69134 36372 69186
rect 36204 69132 36372 69134
rect 36204 68516 36260 69132
rect 37884 68740 37940 70702
rect 37884 68674 37940 68684
rect 36204 68450 36260 68460
rect 38108 60228 38164 73164
rect 38220 73154 38276 73164
rect 38668 73220 38724 73230
rect 38780 73220 38836 73230
rect 38668 73218 38780 73220
rect 38668 73166 38670 73218
rect 38722 73166 38780 73218
rect 38668 73164 38780 73166
rect 38668 73154 38724 73164
rect 38332 72548 38388 72558
rect 38332 72454 38388 72492
rect 38780 72548 38836 73164
rect 38780 72454 38836 72492
rect 39116 73218 39172 73230
rect 39116 73166 39118 73218
rect 39170 73166 39172 73218
rect 38668 72212 38724 72222
rect 38220 71652 38276 71662
rect 38220 71650 38388 71652
rect 38220 71598 38222 71650
rect 38274 71598 38388 71650
rect 38220 71596 38388 71598
rect 38220 71586 38276 71596
rect 38332 71538 38388 71596
rect 38332 71486 38334 71538
rect 38386 71486 38388 71538
rect 38332 70754 38388 71486
rect 38332 70702 38334 70754
rect 38386 70702 38388 70754
rect 38332 63812 38388 70702
rect 38332 63746 38388 63756
rect 38108 60162 38164 60172
rect 38668 58212 38724 72156
rect 39116 66836 39172 73166
rect 39228 73220 39284 73838
rect 39228 73154 39284 73164
rect 39564 73890 40180 73892
rect 39564 73838 39678 73890
rect 39730 73838 40126 73890
rect 40178 73838 40180 73890
rect 39564 73836 40180 73838
rect 39564 73220 39620 73836
rect 39676 73826 39732 73836
rect 40124 73826 40180 73836
rect 39564 73126 39620 73164
rect 40796 68852 40852 74734
rect 41356 72100 41412 74956
rect 41468 74788 41524 74798
rect 41468 74694 41524 74732
rect 41356 72034 41412 72044
rect 41916 71764 41972 75406
rect 42364 73780 42420 76302
rect 42364 73714 42420 73724
rect 46620 76354 46676 76366
rect 46620 76302 46622 76354
rect 46674 76302 46676 76354
rect 46620 72436 46676 76302
rect 46620 72370 46676 72380
rect 41916 71698 41972 71708
rect 40796 68786 40852 68796
rect 39116 66770 39172 66780
rect 38668 57652 38724 58156
rect 40348 66388 40404 66398
rect 38668 57586 38724 57596
rect 40012 57652 40068 57662
rect 36092 51986 36148 51996
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 32620 5236 32676 41916
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34300 5796 34356 5806
rect 34300 5794 34468 5796
rect 34300 5742 34302 5794
rect 34354 5742 34468 5794
rect 34300 5740 34468 5742
rect 34300 5730 34356 5740
rect 33068 5236 33124 5246
rect 32620 5234 33124 5236
rect 32620 5182 32622 5234
rect 32674 5182 33070 5234
rect 33122 5182 33124 5234
rect 32620 5180 33124 5182
rect 32620 5170 32676 5180
rect 33068 5170 33124 5180
rect 34300 5236 34356 5246
rect 34300 5142 34356 5180
rect 27244 4562 27860 4564
rect 27244 4510 27246 4562
rect 27298 4510 27860 4562
rect 27244 4508 27860 4510
rect 27244 4498 27300 4508
rect 27804 4338 27860 4508
rect 27804 4286 27806 4338
rect 27858 4286 27860 4338
rect 27804 4274 27860 4286
rect 28028 5124 28084 5134
rect 28028 4338 28084 5068
rect 32060 5124 32116 5134
rect 32060 5030 32116 5068
rect 33292 5124 33348 5134
rect 33292 5030 33348 5068
rect 34412 5124 34468 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34748 5236 34804 5246
rect 34748 5142 34804 5180
rect 40012 5236 40068 57596
rect 40348 54740 40404 66332
rect 40348 53844 40404 54684
rect 47852 59332 47908 59342
rect 40348 53778 40404 53788
rect 41244 53844 41300 53854
rect 40460 5236 40516 5246
rect 40012 5234 40516 5236
rect 40012 5182 40014 5234
rect 40066 5182 40462 5234
rect 40514 5182 40516 5234
rect 40012 5180 40516 5182
rect 40012 5170 40068 5180
rect 40460 5170 40516 5180
rect 34412 5058 34468 5068
rect 34972 5124 35028 5134
rect 34972 5030 35028 5068
rect 39452 5124 39508 5134
rect 39452 5030 39508 5068
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 33628 4900 33684 4910
rect 33628 4898 34244 4900
rect 33628 4846 33630 4898
rect 33682 4846 34244 4898
rect 33628 4844 34244 4846
rect 33628 4834 33684 4844
rect 29596 4452 29652 4462
rect 29596 4358 29652 4396
rect 30716 4452 30772 4462
rect 34188 4452 34244 4844
rect 35308 4898 35364 4910
rect 35308 4846 35310 4898
rect 35362 4846 35364 4898
rect 34300 4452 34356 4462
rect 34188 4450 34356 4452
rect 34188 4398 34302 4450
rect 34354 4398 34356 4450
rect 34188 4396 34356 4398
rect 28028 4286 28030 4338
rect 28082 4286 28084 4338
rect 28028 4274 28084 4286
rect 28364 4340 28420 4350
rect 28364 4246 28420 4284
rect 29260 4340 29316 4350
rect 29260 4246 29316 4284
rect 26684 3668 26740 3678
rect 26684 3574 26740 3612
rect 30492 3668 30548 3678
rect 26012 3502 26014 3554
rect 26066 3502 26068 3554
rect 26012 3490 26068 3502
rect 30492 800 30548 3612
rect 30716 3554 30772 4396
rect 34300 4386 34356 4396
rect 34636 4450 34692 4462
rect 34636 4398 34638 4450
rect 34690 4398 34692 4450
rect 31388 3668 31444 3678
rect 31388 3574 31444 3612
rect 30716 3502 30718 3554
rect 30770 3502 30772 3554
rect 30716 3490 30772 3502
rect 34636 3556 34692 4398
rect 35308 4452 35364 4846
rect 41020 4898 41076 4910
rect 41020 4846 41022 4898
rect 41074 4846 41076 4898
rect 35308 4386 35364 4396
rect 38332 4452 38388 4462
rect 38332 4358 38388 4396
rect 38668 4450 38724 4462
rect 38668 4398 38670 4450
rect 38722 4398 38724 4450
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35196 3668 35252 3678
rect 35084 3556 35140 3566
rect 34636 3554 35140 3556
rect 34636 3502 35086 3554
rect 35138 3502 35140 3554
rect 34636 3500 35140 3502
rect 35084 3490 35140 3500
rect 35196 800 35252 3612
rect 35756 3668 35812 3678
rect 35756 3574 35812 3612
rect 38668 3556 38724 4398
rect 41020 4452 41076 4846
rect 41020 4386 41076 4396
rect 38668 3490 38724 3500
rect 39900 3668 39956 3678
rect 39900 800 39956 3612
rect 41020 3556 41076 3566
rect 41020 3462 41076 3500
rect 41244 3556 41300 53788
rect 46844 5348 46900 5358
rect 46844 5234 46900 5292
rect 46844 5182 46846 5234
rect 46898 5182 46900 5234
rect 46844 5170 46900 5182
rect 47740 5348 47796 5358
rect 47740 5234 47796 5292
rect 47740 5182 47742 5234
rect 47794 5182 47796 5234
rect 47740 5170 47796 5182
rect 47180 5124 47236 5134
rect 47180 5030 47236 5068
rect 47852 4564 47908 59276
rect 48860 50372 48916 77980
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50876 76580 50932 79200
rect 50876 76514 50932 76524
rect 51548 76580 51604 76590
rect 51548 76486 51604 76524
rect 52668 76580 52724 76590
rect 52668 76486 52724 76524
rect 50540 76356 50596 76366
rect 50428 76354 50596 76356
rect 50428 76302 50542 76354
rect 50594 76302 50596 76354
rect 50428 76300 50596 76302
rect 50428 71876 50484 76300
rect 50540 76290 50596 76300
rect 55020 75796 55076 75806
rect 55244 75796 55300 79200
rect 59612 76692 59668 79200
rect 59948 76692 60004 76702
rect 59612 76690 60004 76692
rect 59612 76638 59950 76690
rect 60002 76638 60004 76690
rect 59612 76636 60004 76638
rect 59948 76580 60004 76636
rect 63868 76692 63924 76702
rect 63980 76692 64036 79200
rect 63868 76690 64036 76692
rect 63868 76638 63870 76690
rect 63922 76638 64036 76690
rect 63868 76636 64036 76638
rect 63868 76626 63924 76636
rect 59948 76514 60004 76524
rect 61628 76580 61684 76590
rect 61628 76486 61684 76524
rect 63980 76580 64036 76636
rect 67788 76804 67844 76814
rect 67788 76690 67844 76748
rect 68348 76804 68404 79200
rect 68348 76738 68404 76748
rect 69580 76804 69636 76814
rect 67788 76638 67790 76690
rect 67842 76638 67844 76690
rect 67788 76626 67844 76638
rect 63980 76514 64036 76524
rect 65548 76580 65604 76590
rect 65548 76486 65604 76524
rect 69580 76578 69636 76748
rect 72492 76692 72548 76702
rect 72716 76692 72772 79200
rect 74956 77364 75012 77374
rect 72492 76690 72772 76692
rect 72492 76638 72494 76690
rect 72546 76638 72772 76690
rect 72492 76636 72772 76638
rect 72492 76626 72548 76636
rect 69580 76526 69582 76578
rect 69634 76526 69636 76578
rect 69580 76514 69636 76526
rect 72716 76580 72772 76636
rect 72716 76514 72772 76524
rect 72940 76692 72996 76702
rect 60620 76354 60676 76366
rect 60620 76302 60622 76354
rect 60674 76302 60676 76354
rect 55468 75796 55524 75806
rect 55020 75794 55300 75796
rect 55020 75742 55022 75794
rect 55074 75742 55300 75794
rect 55020 75740 55300 75742
rect 55020 75730 55076 75740
rect 55244 75572 55300 75740
rect 55244 75506 55300 75516
rect 55356 75794 55524 75796
rect 55356 75742 55470 75794
rect 55522 75742 55524 75794
rect 55356 75740 55524 75742
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 55356 72884 55412 75740
rect 55468 75730 55524 75740
rect 56476 75572 56532 75582
rect 56476 75478 56532 75516
rect 60620 74676 60676 76302
rect 60620 74610 60676 74620
rect 64540 76354 64596 76366
rect 64540 76302 64542 76354
rect 64594 76302 64596 76354
rect 64540 74116 64596 76302
rect 68572 76354 68628 76366
rect 68572 76302 68574 76354
rect 68626 76302 68628 76354
rect 68572 76244 68628 76302
rect 72940 76354 72996 76636
rect 73948 76580 74004 76590
rect 73948 76486 74004 76524
rect 72940 76302 72942 76354
rect 72994 76302 72996 76354
rect 72940 76290 72996 76302
rect 68572 76178 68628 76188
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 74956 75794 75012 77308
rect 74956 75742 74958 75794
rect 75010 75742 75012 75794
rect 74956 75730 75012 75742
rect 77084 75796 77140 79200
rect 77196 75796 77252 75806
rect 77084 75794 77252 75796
rect 77084 75742 77198 75794
rect 77250 75742 77252 75794
rect 77084 75740 77252 75742
rect 76300 75572 76356 75582
rect 77084 75572 77140 75740
rect 77196 75730 77252 75740
rect 76300 75570 77140 75572
rect 76300 75518 76302 75570
rect 76354 75518 77140 75570
rect 76300 75516 77140 75518
rect 76300 75506 76356 75516
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 64540 74050 64596 74060
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 55356 72818 55412 72828
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50428 71810 50484 71820
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 77308 55076 77364 55086
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 48860 49812 48916 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 48860 49746 48916 49756
rect 49532 49812 49588 49822
rect 49532 6132 49588 49756
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49532 6066 49588 6076
rect 51212 6132 51268 6142
rect 51212 6038 51268 6076
rect 52220 6132 52276 6142
rect 52220 5906 52276 6076
rect 52220 5854 52222 5906
rect 52274 5854 52276 5906
rect 52220 5842 52276 5854
rect 52892 5908 52948 5918
rect 51772 5794 51828 5806
rect 51772 5742 51774 5794
rect 51826 5742 51828 5794
rect 47964 5124 48020 5134
rect 47964 5030 48020 5068
rect 51212 5124 51268 5134
rect 47852 4498 47908 4508
rect 48300 4898 48356 4910
rect 48300 4846 48302 4898
rect 48354 4846 48356 4898
rect 43484 4452 43540 4462
rect 43484 4358 43540 4396
rect 43820 4450 43876 4462
rect 43820 4398 43822 4450
rect 43874 4398 43876 4450
rect 41692 3668 41748 3678
rect 41692 3574 41748 3612
rect 43820 3556 43876 4398
rect 48300 4452 48356 4846
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50764 4564 50820 4574
rect 50764 4470 50820 4508
rect 51212 4562 51268 5068
rect 51772 5124 51828 5742
rect 52444 5682 52500 5694
rect 52444 5630 52446 5682
rect 52498 5630 52500 5682
rect 51772 5058 51828 5068
rect 51996 5124 52052 5134
rect 51212 4510 51214 4562
rect 51266 4510 51268 4562
rect 51212 4498 51268 4510
rect 51772 4564 51828 4574
rect 48300 4386 48356 4396
rect 49532 4452 49588 4462
rect 49532 4358 49588 4396
rect 49868 4452 49924 4462
rect 49868 4358 49924 4396
rect 50540 4452 50596 4462
rect 45612 3666 45668 3678
rect 45612 3614 45614 3666
rect 45666 3614 45668 3666
rect 44940 3556 44996 3566
rect 43820 3554 44996 3556
rect 43820 3502 44942 3554
rect 44994 3502 44996 3554
rect 43820 3500 44996 3502
rect 41244 3490 41300 3500
rect 44940 3490 44996 3500
rect 45612 3444 45668 3614
rect 50540 3554 50596 4396
rect 51772 4338 51828 4508
rect 51772 4286 51774 4338
rect 51826 4286 51828 4338
rect 51772 4274 51828 4286
rect 51996 4340 52052 5068
rect 52332 5124 52388 5134
rect 52444 5124 52500 5630
rect 52388 5068 52500 5124
rect 52780 5682 52836 5694
rect 52780 5630 52782 5682
rect 52834 5630 52836 5682
rect 52332 5030 52388 5068
rect 52780 4452 52836 5630
rect 52780 4386 52836 4396
rect 51996 4338 52164 4340
rect 51996 4286 51998 4338
rect 52050 4286 52164 4338
rect 51996 4284 52164 4286
rect 51996 4274 52052 4284
rect 52108 3666 52164 4284
rect 52892 4338 52948 5852
rect 53340 5908 53396 5918
rect 53340 5234 53396 5852
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 53340 5182 53342 5234
rect 53394 5182 53396 5234
rect 53340 5170 53396 5182
rect 52892 4286 52894 4338
rect 52946 4286 52948 4338
rect 52892 4274 52948 4286
rect 53004 5124 53060 5134
rect 53004 4340 53060 5068
rect 54348 4450 54404 4462
rect 54348 4398 54350 4450
rect 54402 4398 54404 4450
rect 53116 4340 53172 4350
rect 53004 4338 53172 4340
rect 53004 4286 53118 4338
rect 53170 4286 53172 4338
rect 53004 4284 53172 4286
rect 52332 4228 52388 4238
rect 52332 4134 52388 4172
rect 53004 3778 53060 4284
rect 53116 4274 53172 4284
rect 53452 4340 53508 4350
rect 53452 4246 53508 4284
rect 54012 4340 54068 4350
rect 54012 4246 54068 4284
rect 53004 3726 53006 3778
rect 53058 3726 53060 3778
rect 53004 3714 53060 3726
rect 52108 3614 52110 3666
rect 52162 3614 52164 3666
rect 52108 3602 52164 3614
rect 54012 3668 54068 3678
rect 50540 3502 50542 3554
rect 50594 3502 50596 3554
rect 50540 3490 50596 3502
rect 51660 3556 51716 3566
rect 51660 3462 51716 3500
rect 52780 3556 52836 3566
rect 52780 3462 52836 3500
rect 53340 3556 53396 3566
rect 53340 3462 53396 3500
rect 49644 3444 49700 3454
rect 45612 3378 45668 3388
rect 49308 3442 49700 3444
rect 49308 3390 49646 3442
rect 49698 3390 49700 3442
rect 49308 3388 49700 3390
rect 44604 3332 44660 3342
rect 44604 800 44660 3276
rect 49308 800 49364 3388
rect 49644 3378 49700 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 54012 800 54068 3612
rect 54348 3554 54404 4398
rect 54908 4452 54964 4462
rect 54908 4358 54964 4396
rect 55244 4452 55300 4462
rect 55244 4358 55300 4396
rect 58268 4452 58324 4462
rect 58268 4358 58324 4396
rect 64540 4452 64596 4462
rect 57932 4338 57988 4350
rect 57932 4286 57934 4338
rect 57986 4286 57988 4338
rect 57932 4228 57988 4286
rect 57932 4162 57988 4172
rect 58604 4340 58660 4350
rect 54908 3668 54964 3678
rect 54908 3574 54964 3612
rect 54348 3502 54350 3554
rect 54402 3502 54404 3554
rect 54348 3490 54404 3502
rect 58604 3554 58660 4284
rect 58604 3502 58606 3554
rect 58658 3502 58660 3554
rect 58604 3490 58660 3502
rect 58716 3668 58772 3678
rect 58716 800 58772 3612
rect 59276 3668 59332 3678
rect 59276 3574 59332 3612
rect 63420 3668 63476 3678
rect 63420 800 63476 3612
rect 64540 3554 64596 4396
rect 66220 4452 66276 4462
rect 66220 4358 66276 4396
rect 68460 4452 68516 4462
rect 65324 4340 65380 4350
rect 65324 4226 65380 4284
rect 65884 4340 65940 4350
rect 65884 4246 65940 4284
rect 65324 4174 65326 4226
rect 65378 4174 65380 4226
rect 65212 3668 65268 3678
rect 65212 3574 65268 3612
rect 64540 3502 64542 3554
rect 64594 3502 64596 3554
rect 64540 3490 64596 3502
rect 65324 3556 65380 4174
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 65324 3490 65380 3500
rect 68124 3668 68180 3678
rect 68124 800 68180 3612
rect 68460 3554 68516 4396
rect 74396 4340 74452 4350
rect 74396 4246 74452 4284
rect 75180 4340 75236 4350
rect 75180 4246 75236 4284
rect 76076 4228 76132 4238
rect 76076 4134 76132 4172
rect 69132 3668 69188 3678
rect 69132 3574 69188 3612
rect 72828 3668 72884 3678
rect 68460 3502 68462 3554
rect 68514 3502 68516 3554
rect 68460 3490 68516 3502
rect 72604 3556 72660 3566
rect 72604 3462 72660 3500
rect 72828 800 72884 3612
rect 73724 3668 73780 3678
rect 73724 3574 73780 3612
rect 73276 3556 73332 3566
rect 73276 3462 73332 3500
rect 77308 3556 77364 55020
rect 77420 36260 77476 36270
rect 77420 4340 77476 36204
rect 77420 4274 77476 4284
rect 77308 3490 77364 3500
rect 77532 4228 77588 4238
rect 77532 800 77588 4172
rect 2240 0 2352 800
rect 6944 0 7056 800
rect 11648 0 11760 800
rect 16352 0 16464 800
rect 21056 0 21168 800
rect 25760 0 25872 800
rect 30464 0 30576 800
rect 35168 0 35280 800
rect 39872 0 39984 800
rect 44576 0 44688 800
rect 49280 0 49392 800
rect 53984 0 54096 800
rect 58688 0 58800 800
rect 63392 0 63504 800
rect 68096 0 68208 800
rect 72800 0 72912 800
rect 77504 0 77616 800
<< via2 >>
rect 2044 78764 2100 78820
rect 2156 77308 2212 77364
rect 2044 76412 2100 76468
rect 2044 75906 2100 75908
rect 2044 75854 2046 75906
rect 2046 75854 2098 75906
rect 2098 75854 2100 75906
rect 2044 75852 2100 75854
rect 2044 75404 2100 75460
rect 1596 74620 1652 74676
rect 1708 70588 1764 70644
rect 1932 73554 1988 73556
rect 1932 73502 1934 73554
rect 1934 73502 1986 73554
rect 1986 73502 1988 73554
rect 1932 73500 1988 73502
rect 2044 72658 2100 72660
rect 2044 72606 2046 72658
rect 2046 72606 2098 72658
rect 2098 72606 2100 72658
rect 2044 72604 2100 72606
rect 1932 72156 1988 72212
rect 2380 78988 2436 79044
rect 3052 79884 3108 79940
rect 2940 78540 2996 78596
rect 2716 77868 2772 77924
rect 2492 77756 2548 77812
rect 2604 75516 2660 75572
rect 2380 74284 2436 74340
rect 2828 75458 2884 75460
rect 2828 75406 2830 75458
rect 2830 75406 2882 75458
rect 2882 75406 2884 75458
rect 2828 75404 2884 75406
rect 2828 74674 2884 74676
rect 2828 74622 2830 74674
rect 2830 74622 2882 74674
rect 2882 74622 2884 74674
rect 2828 74620 2884 74622
rect 2828 74172 2884 74228
rect 2380 71986 2436 71988
rect 2380 71934 2382 71986
rect 2382 71934 2434 71986
rect 2434 71934 2436 71986
rect 2380 71932 2436 71934
rect 2268 70812 2324 70868
rect 2380 70588 2436 70644
rect 1932 69522 1988 69524
rect 1932 69470 1934 69522
rect 1934 69470 1986 69522
rect 1986 69470 1988 69522
rect 1932 69468 1988 69470
rect 2268 70364 2324 70420
rect 4956 79436 5012 79492
rect 4508 79100 4564 79156
rect 4172 78988 4228 79044
rect 3836 78652 3892 78708
rect 3388 78316 3444 78372
rect 3276 76748 3332 76804
rect 3500 76578 3556 76580
rect 3500 76526 3502 76578
rect 3502 76526 3554 76578
rect 3554 76526 3556 76578
rect 3500 76524 3556 76526
rect 3388 75964 3444 76020
rect 3500 76300 3556 76356
rect 3612 76188 3668 76244
rect 2828 73218 2884 73220
rect 2828 73166 2830 73218
rect 2830 73166 2882 73218
rect 2882 73166 2884 73218
rect 2828 73164 2884 73166
rect 2828 71650 2884 71652
rect 2828 71598 2830 71650
rect 2830 71598 2882 71650
rect 2882 71598 2884 71650
rect 2828 71596 2884 71598
rect 2380 70082 2436 70084
rect 2380 70030 2382 70082
rect 2382 70030 2434 70082
rect 2434 70030 2436 70082
rect 2380 70028 2436 70030
rect 2156 69244 2212 69300
rect 2044 68626 2100 68628
rect 2044 68574 2046 68626
rect 2046 68574 2098 68626
rect 2098 68574 2100 68626
rect 2044 68572 2100 68574
rect 1932 68012 1988 68068
rect 1932 67618 1988 67620
rect 1932 67566 1934 67618
rect 1934 67566 1986 67618
rect 1986 67566 1988 67618
rect 1932 67564 1988 67566
rect 2044 67452 2100 67508
rect 1932 65884 1988 65940
rect 1932 65548 1988 65604
rect 2380 68796 2436 68852
rect 2492 69132 2548 69188
rect 2380 67340 2436 67396
rect 2604 67116 2660 67172
rect 2828 69020 2884 69076
rect 3052 69916 3108 69972
rect 3612 75964 3668 76020
rect 3724 75740 3780 75796
rect 3724 75516 3780 75572
rect 4060 77420 4116 77476
rect 3948 76636 4004 76692
rect 4396 76466 4452 76468
rect 4396 76414 4398 76466
rect 4398 76414 4450 76466
rect 4450 76414 4452 76466
rect 4396 76412 4452 76414
rect 4844 78428 4900 78484
rect 4620 77532 4676 77588
rect 4732 77308 4788 77364
rect 4508 76300 4564 76356
rect 4620 76242 4676 76244
rect 4620 76190 4622 76242
rect 4622 76190 4674 76242
rect 4674 76190 4676 76242
rect 4620 76188 4676 76190
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 3948 75516 4004 75572
rect 4508 75682 4564 75684
rect 4508 75630 4510 75682
rect 4510 75630 4562 75682
rect 4562 75630 4564 75682
rect 4508 75628 4564 75630
rect 4396 75516 4452 75572
rect 3836 75404 3892 75460
rect 4732 75570 4788 75572
rect 4732 75518 4734 75570
rect 4734 75518 4786 75570
rect 4786 75518 4788 75570
rect 4732 75516 4788 75518
rect 3500 74002 3556 74004
rect 3500 73950 3502 74002
rect 3502 73950 3554 74002
rect 3554 73950 3556 74002
rect 3500 73948 3556 73950
rect 3388 73500 3444 73556
rect 3276 72380 3332 72436
rect 4060 74956 4116 75012
rect 3948 74002 4004 74004
rect 3948 73950 3950 74002
rect 3950 73950 4002 74002
rect 4002 73950 4004 74002
rect 3948 73948 4004 73950
rect 3836 73836 3892 73892
rect 3724 73218 3780 73220
rect 3724 73166 3726 73218
rect 3726 73166 3778 73218
rect 3778 73166 3780 73218
rect 3724 73164 3780 73166
rect 4172 74732 4228 74788
rect 4508 74732 4564 74788
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 10892 79548 10948 79604
rect 8316 79324 8372 79380
rect 4956 77308 5012 77364
rect 5852 78876 5908 78932
rect 7084 77698 7140 77700
rect 7084 77646 7086 77698
rect 7086 77646 7138 77698
rect 7138 77646 7140 77698
rect 7084 77644 7140 77646
rect 6636 76748 6692 76804
rect 6300 76466 6356 76468
rect 6300 76414 6302 76466
rect 6302 76414 6354 76466
rect 6354 76414 6356 76466
rect 6300 76412 6356 76414
rect 7644 78204 7700 78260
rect 6636 76300 6692 76356
rect 5628 76188 5684 76244
rect 5404 75852 5460 75908
rect 4956 74844 5012 74900
rect 5180 74956 5236 75012
rect 4956 74284 5012 74340
rect 4396 74114 4452 74116
rect 4396 74062 4398 74114
rect 4398 74062 4450 74114
rect 4450 74062 4452 74114
rect 4396 74060 4452 74062
rect 4732 74114 4788 74116
rect 4732 74062 4734 74114
rect 4734 74062 4786 74114
rect 4786 74062 4788 74114
rect 4732 74060 4788 74062
rect 4844 73724 4900 73780
rect 4508 73052 4564 73108
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4284 72716 4340 72772
rect 3724 72604 3780 72660
rect 3388 71762 3444 71764
rect 3388 71710 3390 71762
rect 3390 71710 3442 71762
rect 3442 71710 3444 71762
rect 3388 71708 3444 71710
rect 3388 71484 3444 71540
rect 5292 74844 5348 74900
rect 5292 74060 5348 74116
rect 5180 73330 5236 73332
rect 5180 73278 5182 73330
rect 5182 73278 5234 73330
rect 5234 73278 5236 73330
rect 5180 73276 5236 73278
rect 3836 72546 3892 72548
rect 3836 72494 3838 72546
rect 3838 72494 3890 72546
rect 3890 72494 3892 72546
rect 3836 72492 3892 72494
rect 3164 69522 3220 69524
rect 3164 69470 3166 69522
rect 3166 69470 3218 69522
rect 3218 69470 3220 69522
rect 3164 69468 3220 69470
rect 2940 68684 2996 68740
rect 2828 67842 2884 67844
rect 2828 67790 2830 67842
rect 2830 67790 2882 67842
rect 2882 67790 2884 67842
rect 2828 67788 2884 67790
rect 2268 65490 2324 65492
rect 2268 65438 2270 65490
rect 2270 65438 2322 65490
rect 2322 65438 2324 65490
rect 2268 65436 2324 65438
rect 2380 64818 2436 64820
rect 2380 64766 2382 64818
rect 2382 64766 2434 64818
rect 2434 64766 2436 64818
rect 2380 64764 2436 64766
rect 2156 64092 2212 64148
rect 2268 64652 2324 64708
rect 1820 63980 1876 64036
rect 1932 63756 1988 63812
rect 2380 64204 2436 64260
rect 2380 63922 2436 63924
rect 2380 63870 2382 63922
rect 2382 63870 2434 63922
rect 2434 63870 2436 63922
rect 2380 63868 2436 63870
rect 2716 66444 2772 66500
rect 2604 66386 2660 66388
rect 2604 66334 2606 66386
rect 2606 66334 2658 66386
rect 2658 66334 2660 66386
rect 2604 66332 2660 66334
rect 2716 65100 2772 65156
rect 2492 63532 2548 63588
rect 2940 66892 2996 66948
rect 2828 64764 2884 64820
rect 2940 66444 2996 66500
rect 2828 64594 2884 64596
rect 2828 64542 2830 64594
rect 2830 64542 2882 64594
rect 2882 64542 2884 64594
rect 2828 64540 2884 64542
rect 2380 63138 2436 63140
rect 2380 63086 2382 63138
rect 2382 63086 2434 63138
rect 2434 63086 2436 63138
rect 2380 63084 2436 63086
rect 3388 68684 3444 68740
rect 3164 68012 3220 68068
rect 3388 67900 3444 67956
rect 3276 67730 3332 67732
rect 3276 67678 3278 67730
rect 3278 67678 3330 67730
rect 3330 67678 3332 67730
rect 3276 67676 3332 67678
rect 3164 67340 3220 67396
rect 3164 67170 3220 67172
rect 3164 67118 3166 67170
rect 3166 67118 3218 67170
rect 3218 67118 3220 67170
rect 3164 67116 3220 67118
rect 3724 71820 3780 71876
rect 3836 71762 3892 71764
rect 3836 71710 3838 71762
rect 3838 71710 3890 71762
rect 3890 71710 3892 71762
rect 3836 71708 3892 71710
rect 4956 73164 5012 73220
rect 4844 72156 4900 72212
rect 4732 71596 4788 71652
rect 4508 71484 4564 71540
rect 3948 71090 4004 71092
rect 3948 71038 3950 71090
rect 3950 71038 4002 71090
rect 4002 71038 4004 71090
rect 3948 71036 4004 71038
rect 3836 70194 3892 70196
rect 3836 70142 3838 70194
rect 3838 70142 3890 70194
rect 3890 70142 3892 70194
rect 3836 70140 3892 70142
rect 3724 69410 3780 69412
rect 3724 69358 3726 69410
rect 3726 69358 3778 69410
rect 3778 69358 3780 69410
rect 3724 69356 3780 69358
rect 3612 68684 3668 68740
rect 3724 68796 3780 68852
rect 3836 68684 3892 68740
rect 3724 68124 3780 68180
rect 3836 67228 3892 67284
rect 3724 67116 3780 67172
rect 3164 66444 3220 66500
rect 3052 65660 3108 65716
rect 3052 65100 3108 65156
rect 3724 66892 3780 66948
rect 3164 64876 3220 64932
rect 3164 64706 3220 64708
rect 3164 64654 3166 64706
rect 3166 64654 3218 64706
rect 3218 64654 3220 64706
rect 3164 64652 3220 64654
rect 3164 63810 3220 63812
rect 3164 63758 3166 63810
rect 3166 63758 3218 63810
rect 3218 63758 3220 63810
rect 3164 63756 3220 63758
rect 2716 63420 2772 63476
rect 2716 62748 2772 62804
rect 2604 62636 2660 62692
rect 3164 63532 3220 63588
rect 3388 64428 3444 64484
rect 3164 62748 3220 62804
rect 3276 62636 3332 62692
rect 1932 61346 1988 61348
rect 1932 61294 1934 61346
rect 1934 61294 1986 61346
rect 1986 61294 1988 61346
rect 1932 61292 1988 61294
rect 1932 61010 1988 61012
rect 1932 60958 1934 61010
rect 1934 60958 1986 61010
rect 1986 60958 1988 61010
rect 1932 60956 1988 60958
rect 1596 60060 1652 60116
rect 2828 62300 2884 62356
rect 2492 61740 2548 61796
rect 2604 62188 2660 62244
rect 2380 61682 2436 61684
rect 2380 61630 2382 61682
rect 2382 61630 2434 61682
rect 2434 61630 2436 61682
rect 2380 61628 2436 61630
rect 3052 62300 3108 62356
rect 2716 61516 2772 61572
rect 2604 60172 2660 60228
rect 2492 59836 2548 59892
rect 2828 62132 2884 62188
rect 3612 64706 3668 64708
rect 3612 64654 3614 64706
rect 3614 64654 3666 64706
rect 3666 64654 3668 64706
rect 3612 64652 3668 64654
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 4172 71148 4228 71204
rect 4844 71148 4900 71204
rect 4620 71090 4676 71092
rect 4620 71038 4622 71090
rect 4622 71038 4674 71090
rect 4674 71038 4676 71090
rect 4620 71036 4676 71038
rect 4396 70978 4452 70980
rect 4396 70926 4398 70978
rect 4398 70926 4450 70978
rect 4450 70926 4452 70978
rect 4396 70924 4452 70926
rect 5516 73106 5572 73108
rect 5516 73054 5518 73106
rect 5518 73054 5570 73106
rect 5570 73054 5572 73106
rect 5516 73052 5572 73054
rect 5068 71820 5124 71876
rect 4956 71036 5012 71092
rect 4844 70924 4900 70980
rect 4396 70476 4452 70532
rect 4956 70754 5012 70756
rect 4956 70702 4958 70754
rect 4958 70702 5010 70754
rect 5010 70702 5012 70754
rect 4956 70700 5012 70702
rect 5292 72492 5348 72548
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 4508 69522 4564 69524
rect 4508 69470 4510 69522
rect 4510 69470 4562 69522
rect 4562 69470 4564 69522
rect 4508 69468 4564 69470
rect 4284 69244 4340 69300
rect 4844 69132 4900 69188
rect 4396 68738 4452 68740
rect 4396 68686 4398 68738
rect 4398 68686 4450 68738
rect 4450 68686 4452 68738
rect 4396 68684 4452 68686
rect 4844 68572 4900 68628
rect 5180 70028 5236 70084
rect 5068 69692 5124 69748
rect 4284 68236 4340 68292
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 4844 68124 4900 68180
rect 5068 69132 5124 69188
rect 4620 67842 4676 67844
rect 4620 67790 4622 67842
rect 4622 67790 4674 67842
rect 4674 67790 4676 67842
rect 4620 67788 4676 67790
rect 5404 72044 5460 72100
rect 6300 76188 6356 76244
rect 5964 75852 6020 75908
rect 5740 74172 5796 74228
rect 6076 74620 6132 74676
rect 6188 73500 6244 73556
rect 6748 76076 6804 76132
rect 7308 76412 7364 76468
rect 6412 73890 6468 73892
rect 6412 73838 6414 73890
rect 6414 73838 6466 73890
rect 6466 73838 6468 73890
rect 6412 73836 6468 73838
rect 6188 73330 6244 73332
rect 6188 73278 6190 73330
rect 6190 73278 6242 73330
rect 6242 73278 6244 73330
rect 6188 73276 6244 73278
rect 6412 73330 6468 73332
rect 6412 73278 6414 73330
rect 6414 73278 6466 73330
rect 6466 73278 6468 73330
rect 6412 73276 6468 73278
rect 5740 72044 5796 72100
rect 5852 73052 5908 73108
rect 6300 72770 6356 72772
rect 6300 72718 6302 72770
rect 6302 72718 6354 72770
rect 6354 72718 6356 72770
rect 6300 72716 6356 72718
rect 6188 72492 6244 72548
rect 5740 71874 5796 71876
rect 5740 71822 5742 71874
rect 5742 71822 5794 71874
rect 5794 71822 5796 71874
rect 5740 71820 5796 71822
rect 5404 70700 5460 70756
rect 5516 71484 5572 71540
rect 5068 68572 5124 68628
rect 4284 67116 4340 67172
rect 4172 66946 4228 66948
rect 4172 66894 4174 66946
rect 4174 66894 4226 66946
rect 4226 66894 4228 66946
rect 4172 66892 4228 66894
rect 4060 66386 4116 66388
rect 4060 66334 4062 66386
rect 4062 66334 4114 66386
rect 4114 66334 4116 66386
rect 4060 66332 4116 66334
rect 3836 65436 3892 65492
rect 4060 65490 4116 65492
rect 4060 65438 4062 65490
rect 4062 65438 4114 65490
rect 4114 65438 4116 65490
rect 4060 65436 4116 65438
rect 4060 64482 4116 64484
rect 4060 64430 4062 64482
rect 4062 64430 4114 64482
rect 4114 64430 4116 64482
rect 4060 64428 4116 64430
rect 3612 63980 3668 64036
rect 3948 63980 4004 64036
rect 3724 63922 3780 63924
rect 3724 63870 3726 63922
rect 3726 63870 3778 63922
rect 3778 63870 3780 63922
rect 3724 63868 3780 63870
rect 3500 63420 3556 63476
rect 3164 61740 3220 61796
rect 3164 61180 3220 61236
rect 3276 60956 3332 61012
rect 3052 60114 3108 60116
rect 3052 60062 3054 60114
rect 3054 60062 3106 60114
rect 3106 60062 3108 60114
rect 3052 60060 3108 60062
rect 3612 63308 3668 63364
rect 3724 61740 3780 61796
rect 3612 61346 3668 61348
rect 3612 61294 3614 61346
rect 3614 61294 3666 61346
rect 3666 61294 3668 61346
rect 3612 61292 3668 61294
rect 3724 60732 3780 60788
rect 3052 59276 3108 59332
rect 3388 59388 3444 59444
rect 4508 67116 4564 67172
rect 4956 67116 5012 67172
rect 4620 67058 4676 67060
rect 4620 67006 4622 67058
rect 4622 67006 4674 67058
rect 4674 67006 4676 67058
rect 4620 67004 4676 67006
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 5404 69468 5460 69524
rect 5404 68908 5460 68964
rect 5292 68402 5348 68404
rect 5292 68350 5294 68402
rect 5294 68350 5346 68402
rect 5346 68350 5348 68402
rect 5292 68348 5348 68350
rect 6188 72322 6244 72324
rect 6188 72270 6190 72322
rect 6190 72270 6242 72322
rect 6242 72270 6244 72322
rect 6188 72268 6244 72270
rect 6300 72156 6356 72212
rect 6188 72044 6244 72100
rect 5964 71762 6020 71764
rect 5964 71710 5966 71762
rect 5966 71710 6018 71762
rect 6018 71710 6020 71762
rect 5964 71708 6020 71710
rect 5964 71372 6020 71428
rect 5852 70700 5908 70756
rect 6860 75628 6916 75684
rect 7196 75516 7252 75572
rect 7084 74396 7140 74452
rect 6972 73948 7028 74004
rect 7196 73948 7252 74004
rect 6748 73836 6804 73892
rect 6972 73500 7028 73556
rect 6636 72604 6692 72660
rect 6860 72546 6916 72548
rect 6860 72494 6862 72546
rect 6862 72494 6914 72546
rect 6914 72494 6916 72546
rect 6860 72492 6916 72494
rect 6300 71260 6356 71316
rect 6412 71036 6468 71092
rect 6524 70978 6580 70980
rect 6524 70926 6526 70978
rect 6526 70926 6578 70978
rect 6578 70926 6580 70978
rect 6524 70924 6580 70926
rect 5628 70418 5684 70420
rect 5628 70366 5630 70418
rect 5630 70366 5682 70418
rect 5682 70366 5684 70418
rect 5628 70364 5684 70366
rect 6076 70588 6132 70644
rect 5628 69692 5684 69748
rect 5852 69634 5908 69636
rect 5852 69582 5854 69634
rect 5854 69582 5906 69634
rect 5906 69582 5908 69634
rect 5852 69580 5908 69582
rect 5740 69244 5796 69300
rect 6300 70364 6356 70420
rect 6412 70700 6468 70756
rect 6188 70252 6244 70308
rect 6300 69634 6356 69636
rect 6300 69582 6302 69634
rect 6302 69582 6354 69634
rect 6354 69582 6356 69634
rect 6300 69580 6356 69582
rect 5964 68684 6020 68740
rect 6076 69244 6132 69300
rect 5180 66892 5236 66948
rect 4956 66556 5012 66612
rect 4508 66444 4564 66500
rect 4284 66108 4340 66164
rect 4396 65996 4452 66052
rect 4508 65772 4564 65828
rect 4620 65884 4676 65940
rect 5068 65772 5124 65828
rect 5852 66946 5908 66948
rect 5852 66894 5854 66946
rect 5854 66894 5906 66946
rect 5906 66894 5908 66946
rect 5852 66892 5908 66894
rect 5516 65772 5572 65828
rect 5628 65660 5684 65716
rect 4844 65602 4900 65604
rect 4844 65550 4846 65602
rect 4846 65550 4898 65602
rect 4898 65550 4900 65602
rect 4844 65548 4900 65550
rect 5404 65548 5460 65604
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 4956 64988 5012 65044
rect 4508 64594 4564 64596
rect 4508 64542 4510 64594
rect 4510 64542 4562 64594
rect 4562 64542 4564 64594
rect 4508 64540 4564 64542
rect 4956 64818 5012 64820
rect 4956 64766 4958 64818
rect 4958 64766 5010 64818
rect 5010 64766 5012 64818
rect 4956 64764 5012 64766
rect 5516 65266 5572 65268
rect 5516 65214 5518 65266
rect 5518 65214 5570 65266
rect 5570 65214 5572 65266
rect 5516 65212 5572 65214
rect 5180 64540 5236 64596
rect 4844 64428 4900 64484
rect 5740 65324 5796 65380
rect 5852 65660 5908 65716
rect 5516 64146 5572 64148
rect 5516 64094 5518 64146
rect 5518 64094 5570 64146
rect 5570 64094 5572 64146
rect 5516 64092 5572 64094
rect 4172 63644 4228 63700
rect 4844 63756 4900 63812
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4172 63308 4228 63364
rect 4620 63250 4676 63252
rect 4620 63198 4622 63250
rect 4622 63198 4674 63250
rect 4674 63198 4676 63250
rect 4620 63196 4676 63198
rect 4508 62748 4564 62804
rect 4956 62354 5012 62356
rect 4956 62302 4958 62354
rect 4958 62302 5010 62354
rect 5010 62302 5012 62354
rect 4956 62300 5012 62302
rect 4172 62242 4228 62244
rect 4172 62190 4174 62242
rect 4174 62190 4226 62242
rect 4226 62190 4228 62242
rect 4172 62188 4228 62190
rect 4844 62076 4900 62132
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4172 61628 4228 61684
rect 4060 61570 4116 61572
rect 4060 61518 4062 61570
rect 4062 61518 4114 61570
rect 4114 61518 4116 61570
rect 4060 61516 4116 61518
rect 4508 61682 4564 61684
rect 4508 61630 4510 61682
rect 4510 61630 4562 61682
rect 4562 61630 4564 61682
rect 4508 61628 4564 61630
rect 4396 61180 4452 61236
rect 4060 60620 4116 60676
rect 3724 58604 3780 58660
rect 5852 63196 5908 63252
rect 6300 67452 6356 67508
rect 6076 67116 6132 67172
rect 6076 65660 6132 65716
rect 6748 70588 6804 70644
rect 6748 70418 6804 70420
rect 6748 70366 6750 70418
rect 6750 70366 6802 70418
rect 6802 70366 6804 70418
rect 6748 70364 6804 70366
rect 6636 69692 6692 69748
rect 6524 69132 6580 69188
rect 6636 69244 6692 69300
rect 6188 67228 6244 67284
rect 5964 64764 6020 64820
rect 6524 67564 6580 67620
rect 6636 67116 6692 67172
rect 6524 65660 6580 65716
rect 6300 64764 6356 64820
rect 6300 64540 6356 64596
rect 6860 67452 6916 67508
rect 7084 73052 7140 73108
rect 7196 71762 7252 71764
rect 7196 71710 7198 71762
rect 7198 71710 7250 71762
rect 7250 71710 7252 71762
rect 7196 71708 7252 71710
rect 7196 71484 7252 71540
rect 7532 75404 7588 75460
rect 7532 74674 7588 74676
rect 7532 74622 7534 74674
rect 7534 74622 7586 74674
rect 7586 74622 7588 74674
rect 7532 74620 7588 74622
rect 7980 75740 8036 75796
rect 7756 75010 7812 75012
rect 7756 74958 7758 75010
rect 7758 74958 7810 75010
rect 7810 74958 7812 75010
rect 7756 74956 7812 74958
rect 7644 74114 7700 74116
rect 7644 74062 7646 74114
rect 7646 74062 7698 74114
rect 7698 74062 7700 74114
rect 7644 74060 7700 74062
rect 7420 73724 7476 73780
rect 7644 73612 7700 73668
rect 7980 73948 8036 74004
rect 8204 75794 8260 75796
rect 8204 75742 8206 75794
rect 8206 75742 8258 75794
rect 8258 75742 8260 75794
rect 8204 75740 8260 75742
rect 8204 75292 8260 75348
rect 8204 74060 8260 74116
rect 7868 73500 7924 73556
rect 7420 73052 7476 73108
rect 7420 71596 7476 71652
rect 7308 70924 7364 70980
rect 7308 70476 7364 70532
rect 7420 70588 7476 70644
rect 7308 70082 7364 70084
rect 7308 70030 7310 70082
rect 7310 70030 7362 70082
rect 7362 70030 7364 70082
rect 7308 70028 7364 70030
rect 7532 70082 7588 70084
rect 7532 70030 7534 70082
rect 7534 70030 7586 70082
rect 7586 70030 7588 70082
rect 7532 70028 7588 70030
rect 7196 68348 7252 68404
rect 6748 66556 6804 66612
rect 6860 66162 6916 66164
rect 6860 66110 6862 66162
rect 6862 66110 6914 66162
rect 6914 66110 6916 66162
rect 6860 66108 6916 66110
rect 6636 65324 6692 65380
rect 6748 65100 6804 65156
rect 6860 63922 6916 63924
rect 6860 63870 6862 63922
rect 6862 63870 6914 63922
rect 6914 63870 6916 63922
rect 6860 63868 6916 63870
rect 6300 63756 6356 63812
rect 6636 63196 6692 63252
rect 6300 62860 6356 62916
rect 6412 62578 6468 62580
rect 6412 62526 6414 62578
rect 6414 62526 6466 62578
rect 6466 62526 6468 62578
rect 6412 62524 6468 62526
rect 6076 62076 6132 62132
rect 5852 61740 5908 61796
rect 4956 61180 5012 61236
rect 5964 61516 6020 61572
rect 5292 61068 5348 61124
rect 4172 58940 4228 58996
rect 4956 61010 5012 61012
rect 4956 60958 4958 61010
rect 4958 60958 5010 61010
rect 5010 60958 5012 61010
rect 4956 60956 5012 60958
rect 3388 57820 3444 57876
rect 2940 57708 2996 57764
rect 2828 54460 2884 54516
rect 2716 49980 2772 50036
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4396 59948 4452 60004
rect 4396 59778 4452 59780
rect 4396 59726 4398 59778
rect 4398 59726 4450 59778
rect 4450 59726 4452 59778
rect 4396 59724 4452 59726
rect 4732 59836 4788 59892
rect 4844 59724 4900 59780
rect 4396 59106 4452 59108
rect 4396 59054 4398 59106
rect 4398 59054 4450 59106
rect 4450 59054 4452 59106
rect 4396 59052 4452 59054
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4956 59388 5012 59444
rect 5852 61068 5908 61124
rect 5516 60786 5572 60788
rect 5516 60734 5518 60786
rect 5518 60734 5570 60786
rect 5570 60734 5572 60786
rect 5516 60732 5572 60734
rect 5852 59500 5908 59556
rect 6300 61292 6356 61348
rect 6300 60786 6356 60788
rect 6300 60734 6302 60786
rect 6302 60734 6354 60786
rect 6354 60734 6356 60786
rect 6300 60732 6356 60734
rect 6188 60060 6244 60116
rect 6300 60002 6356 60004
rect 6300 59950 6302 60002
rect 6302 59950 6354 60002
rect 6354 59950 6356 60002
rect 6300 59948 6356 59950
rect 5852 58546 5908 58548
rect 5852 58494 5854 58546
rect 5854 58494 5906 58546
rect 5906 58494 5908 58546
rect 5852 58492 5908 58494
rect 4844 56812 4900 56868
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 6076 58994 6132 58996
rect 6076 58942 6078 58994
rect 6078 58942 6130 58994
rect 6130 58942 6132 58994
rect 6076 58940 6132 58942
rect 6300 58940 6356 58996
rect 6300 58716 6356 58772
rect 6860 63250 6916 63252
rect 6860 63198 6862 63250
rect 6862 63198 6914 63250
rect 6914 63198 6916 63250
rect 6860 63196 6916 63198
rect 7308 67618 7364 67620
rect 7308 67566 7310 67618
rect 7310 67566 7362 67618
rect 7362 67566 7364 67618
rect 7308 67564 7364 67566
rect 7420 67170 7476 67172
rect 7420 67118 7422 67170
rect 7422 67118 7474 67170
rect 7474 67118 7476 67170
rect 7420 67116 7476 67118
rect 7308 66834 7364 66836
rect 7308 66782 7310 66834
rect 7310 66782 7362 66834
rect 7362 66782 7364 66834
rect 7308 66780 7364 66782
rect 7084 65996 7140 66052
rect 7196 66220 7252 66276
rect 7532 66050 7588 66052
rect 7532 65998 7534 66050
rect 7534 65998 7586 66050
rect 7586 65998 7588 66050
rect 7532 65996 7588 65998
rect 7644 65660 7700 65716
rect 7196 64316 7252 64372
rect 7196 63420 7252 63476
rect 7308 63532 7364 63588
rect 7308 63308 7364 63364
rect 7308 62914 7364 62916
rect 7308 62862 7310 62914
rect 7310 62862 7362 62914
rect 7362 62862 7364 62914
rect 7308 62860 7364 62862
rect 7644 64540 7700 64596
rect 7980 72380 8036 72436
rect 7868 72268 7924 72324
rect 8204 72546 8260 72548
rect 8204 72494 8206 72546
rect 8206 72494 8258 72546
rect 8258 72494 8260 72546
rect 8204 72492 8260 72494
rect 8204 72268 8260 72324
rect 7868 71484 7924 71540
rect 7980 71708 8036 71764
rect 7868 69410 7924 69412
rect 7868 69358 7870 69410
rect 7870 69358 7922 69410
rect 7922 69358 7924 69410
rect 7868 69356 7924 69358
rect 8092 70924 8148 70980
rect 8092 70754 8148 70756
rect 8092 70702 8094 70754
rect 8094 70702 8146 70754
rect 8146 70702 8148 70754
rect 8092 70700 8148 70702
rect 8876 79212 8932 79268
rect 8428 77756 8484 77812
rect 8428 76524 8484 76580
rect 9100 77756 9156 77812
rect 8988 75682 9044 75684
rect 8988 75630 8990 75682
rect 8990 75630 9042 75682
rect 9042 75630 9044 75682
rect 8988 75628 9044 75630
rect 8764 75404 8820 75460
rect 8652 74956 8708 75012
rect 8428 74284 8484 74340
rect 8764 74898 8820 74900
rect 8764 74846 8766 74898
rect 8766 74846 8818 74898
rect 8818 74846 8820 74898
rect 8764 74844 8820 74846
rect 8988 74898 9044 74900
rect 8988 74846 8990 74898
rect 8990 74846 9042 74898
rect 9042 74846 9044 74898
rect 8988 74844 9044 74846
rect 8652 74172 8708 74228
rect 8540 73612 8596 73668
rect 8876 73836 8932 73892
rect 8540 73106 8596 73108
rect 8540 73054 8542 73106
rect 8542 73054 8594 73106
rect 8594 73054 8596 73106
rect 8540 73052 8596 73054
rect 8316 70700 8372 70756
rect 8428 72940 8484 72996
rect 8316 70418 8372 70420
rect 8316 70366 8318 70418
rect 8318 70366 8370 70418
rect 8370 70366 8372 70418
rect 8316 70364 8372 70366
rect 8988 73612 9044 73668
rect 9660 77196 9716 77252
rect 10220 77420 10276 77476
rect 9996 76860 10052 76916
rect 10108 75682 10164 75684
rect 10108 75630 10110 75682
rect 10110 75630 10162 75682
rect 10162 75630 10164 75682
rect 10108 75628 10164 75630
rect 9436 73836 9492 73892
rect 8652 72716 8708 72772
rect 8540 71650 8596 71652
rect 8540 71598 8542 71650
rect 8542 71598 8594 71650
rect 8594 71598 8596 71650
rect 8540 71596 8596 71598
rect 8540 70418 8596 70420
rect 8540 70366 8542 70418
rect 8542 70366 8594 70418
rect 8594 70366 8596 70418
rect 8540 70364 8596 70366
rect 8428 70252 8484 70308
rect 8204 70194 8260 70196
rect 8204 70142 8206 70194
rect 8206 70142 8258 70194
rect 8258 70142 8260 70194
rect 8204 70140 8260 70142
rect 8428 70082 8484 70084
rect 8428 70030 8430 70082
rect 8430 70030 8482 70082
rect 8482 70030 8484 70082
rect 8428 70028 8484 70030
rect 8204 69410 8260 69412
rect 8204 69358 8206 69410
rect 8206 69358 8258 69410
rect 8258 69358 8260 69410
rect 8204 69356 8260 69358
rect 8204 68514 8260 68516
rect 8204 68462 8206 68514
rect 8206 68462 8258 68514
rect 8258 68462 8260 68514
rect 8204 68460 8260 68462
rect 8876 71372 8932 71428
rect 8764 70028 8820 70084
rect 8876 68796 8932 68852
rect 8876 68012 8932 68068
rect 9324 73052 9380 73108
rect 9100 72546 9156 72548
rect 9100 72494 9102 72546
rect 9102 72494 9154 72546
rect 9154 72494 9156 72546
rect 9100 72492 9156 72494
rect 9100 71372 9156 71428
rect 9100 70364 9156 70420
rect 9100 69692 9156 69748
rect 9212 69580 9268 69636
rect 8988 67340 9044 67396
rect 8876 67282 8932 67284
rect 8876 67230 8878 67282
rect 8878 67230 8930 67282
rect 8930 67230 8932 67282
rect 8876 67228 8932 67230
rect 8092 66498 8148 66500
rect 8092 66446 8094 66498
rect 8094 66446 8146 66498
rect 8146 66446 8148 66498
rect 8092 66444 8148 66446
rect 8316 66444 8372 66500
rect 7868 66332 7924 66388
rect 7868 64482 7924 64484
rect 7868 64430 7870 64482
rect 7870 64430 7922 64482
rect 7922 64430 7924 64482
rect 7868 64428 7924 64430
rect 6860 61852 6916 61908
rect 6636 61628 6692 61684
rect 6972 61740 7028 61796
rect 6748 61068 6804 61124
rect 6860 61010 6916 61012
rect 6860 60958 6862 61010
rect 6862 60958 6914 61010
rect 6914 60958 6916 61010
rect 6860 60956 6916 60958
rect 7196 61682 7252 61684
rect 7196 61630 7198 61682
rect 7198 61630 7250 61682
rect 7250 61630 7252 61682
rect 7196 61628 7252 61630
rect 7420 62524 7476 62580
rect 7308 61180 7364 61236
rect 7196 60674 7252 60676
rect 7196 60622 7198 60674
rect 7198 60622 7250 60674
rect 7250 60622 7252 60674
rect 7196 60620 7252 60622
rect 7084 59778 7140 59780
rect 7084 59726 7086 59778
rect 7086 59726 7138 59778
rect 7138 59726 7140 59778
rect 7084 59724 7140 59726
rect 7308 59442 7364 59444
rect 7308 59390 7310 59442
rect 7310 59390 7362 59442
rect 7362 59390 7364 59442
rect 7308 59388 7364 59390
rect 6636 58716 6692 58772
rect 6412 56252 6468 56308
rect 6636 58156 6692 58212
rect 7196 58044 7252 58100
rect 7308 57538 7364 57540
rect 7308 57486 7310 57538
rect 7310 57486 7362 57538
rect 7362 57486 7364 57538
rect 7308 57484 7364 57486
rect 6636 51884 6692 51940
rect 8092 65714 8148 65716
rect 8092 65662 8094 65714
rect 8094 65662 8146 65714
rect 8146 65662 8148 65714
rect 8092 65660 8148 65662
rect 8316 65714 8372 65716
rect 8316 65662 8318 65714
rect 8318 65662 8370 65714
rect 8370 65662 8372 65714
rect 8316 65660 8372 65662
rect 8204 65602 8260 65604
rect 8204 65550 8206 65602
rect 8206 65550 8258 65602
rect 8258 65550 8260 65602
rect 8204 65548 8260 65550
rect 8092 64316 8148 64372
rect 8204 64876 8260 64932
rect 7980 63756 8036 63812
rect 7644 63532 7700 63588
rect 7756 63644 7812 63700
rect 7532 61628 7588 61684
rect 7644 62524 7700 62580
rect 7868 63138 7924 63140
rect 7868 63086 7870 63138
rect 7870 63086 7922 63138
rect 7922 63086 7924 63138
rect 7868 63084 7924 63086
rect 8092 62524 8148 62580
rect 8204 63420 8260 63476
rect 8540 65100 8596 65156
rect 8540 64876 8596 64932
rect 8652 66556 8708 66612
rect 8316 63196 8372 63252
rect 8428 63756 8484 63812
rect 8540 63698 8596 63700
rect 8540 63646 8542 63698
rect 8542 63646 8594 63698
rect 8594 63646 8596 63698
rect 8540 63644 8596 63646
rect 8876 66108 8932 66164
rect 8764 65490 8820 65492
rect 8764 65438 8766 65490
rect 8766 65438 8818 65490
rect 8818 65438 8820 65490
rect 8764 65436 8820 65438
rect 8764 65100 8820 65156
rect 8764 64316 8820 64372
rect 8988 66892 9044 66948
rect 9436 72604 9492 72660
rect 9884 74956 9940 75012
rect 9660 74338 9716 74340
rect 9660 74286 9662 74338
rect 9662 74286 9714 74338
rect 9714 74286 9716 74338
rect 9660 74284 9716 74286
rect 9996 74284 10052 74340
rect 10108 74002 10164 74004
rect 10108 73950 10110 74002
rect 10110 73950 10162 74002
rect 10162 73950 10164 74002
rect 10108 73948 10164 73950
rect 9996 73724 10052 73780
rect 10332 74674 10388 74676
rect 10332 74622 10334 74674
rect 10334 74622 10386 74674
rect 10386 74622 10388 74674
rect 10332 74620 10388 74622
rect 10220 73724 10276 73780
rect 10668 76188 10724 76244
rect 14364 79884 14420 79940
rect 10892 75964 10948 76020
rect 11452 77308 11508 77364
rect 10556 75740 10612 75796
rect 10668 75852 10724 75908
rect 10556 74786 10612 74788
rect 10556 74734 10558 74786
rect 10558 74734 10610 74786
rect 10610 74734 10612 74786
rect 10556 74732 10612 74734
rect 10444 73836 10500 73892
rect 10332 73612 10388 73668
rect 10220 73276 10276 73332
rect 10108 73164 10164 73220
rect 9772 71986 9828 71988
rect 9772 71934 9774 71986
rect 9774 71934 9826 71986
rect 9826 71934 9828 71986
rect 9772 71932 9828 71934
rect 9996 71708 10052 71764
rect 9436 69580 9492 69636
rect 9660 69804 9716 69860
rect 10220 71538 10276 71540
rect 10220 71486 10222 71538
rect 10222 71486 10274 71538
rect 10274 71486 10276 71538
rect 10220 71484 10276 71486
rect 10668 73724 10724 73780
rect 10668 73164 10724 73220
rect 10444 72716 10500 72772
rect 11340 75404 11396 75460
rect 12124 77532 12180 77588
rect 12012 76860 12068 76916
rect 11564 76636 11620 76692
rect 11564 76076 11620 76132
rect 11116 74898 11172 74900
rect 11116 74846 11118 74898
rect 11118 74846 11170 74898
rect 11170 74846 11172 74898
rect 11116 74844 11172 74846
rect 11116 74172 11172 74228
rect 11004 74114 11060 74116
rect 11004 74062 11006 74114
rect 11006 74062 11058 74114
rect 11058 74062 11060 74114
rect 11004 74060 11060 74062
rect 10556 72268 10612 72324
rect 9996 70140 10052 70196
rect 9884 69804 9940 69860
rect 9660 69580 9716 69636
rect 9548 69410 9604 69412
rect 9548 69358 9550 69410
rect 9550 69358 9602 69410
rect 9602 69358 9604 69410
rect 9548 69356 9604 69358
rect 9324 68460 9380 68516
rect 9436 68908 9492 68964
rect 9324 68012 9380 68068
rect 9324 66556 9380 66612
rect 9100 66220 9156 66276
rect 8988 64652 9044 64708
rect 8988 64482 9044 64484
rect 8988 64430 8990 64482
rect 8990 64430 9042 64482
rect 9042 64430 9044 64482
rect 8988 64428 9044 64430
rect 9772 69244 9828 69300
rect 9884 69132 9940 69188
rect 10108 68796 10164 68852
rect 9660 68572 9716 68628
rect 10108 68572 10164 68628
rect 9548 67228 9604 67284
rect 9548 66780 9604 66836
rect 9884 67452 9940 67508
rect 9100 64092 9156 64148
rect 9660 65996 9716 66052
rect 8764 63532 8820 63588
rect 8876 63308 8932 63364
rect 8428 62860 8484 62916
rect 8988 62972 9044 63028
rect 8540 62636 8596 62692
rect 8204 62188 8260 62244
rect 8876 62188 8932 62244
rect 7756 61740 7812 61796
rect 8428 61740 8484 61796
rect 7644 61292 7700 61348
rect 7756 60898 7812 60900
rect 7756 60846 7758 60898
rect 7758 60846 7810 60898
rect 7810 60846 7812 60898
rect 7756 60844 7812 60846
rect 7756 60508 7812 60564
rect 8428 61346 8484 61348
rect 8428 61294 8430 61346
rect 8430 61294 8482 61346
rect 8482 61294 8484 61346
rect 8428 61292 8484 61294
rect 8316 61180 8372 61236
rect 7868 60396 7924 60452
rect 8092 60674 8148 60676
rect 8092 60622 8094 60674
rect 8094 60622 8146 60674
rect 8146 60622 8148 60674
rect 8092 60620 8148 60622
rect 7756 60172 7812 60228
rect 8204 60172 8260 60228
rect 8092 59724 8148 59780
rect 7644 59500 7700 59556
rect 7980 59164 8036 59220
rect 7644 58210 7700 58212
rect 7644 58158 7646 58210
rect 7646 58158 7698 58210
rect 7698 58158 7700 58210
rect 7644 58156 7700 58158
rect 7868 57874 7924 57876
rect 7868 57822 7870 57874
rect 7870 57822 7922 57874
rect 7922 57822 7924 57874
rect 7868 57820 7924 57822
rect 7980 56476 8036 56532
rect 8092 57260 8148 57316
rect 8652 61068 8708 61124
rect 8988 60956 9044 61012
rect 8652 60732 8708 60788
rect 8428 60508 8484 60564
rect 8988 60508 9044 60564
rect 8652 60172 8708 60228
rect 9212 63644 9268 63700
rect 9436 65324 9492 65380
rect 10108 68012 10164 68068
rect 10332 70588 10388 70644
rect 10444 70252 10500 70308
rect 11004 72434 11060 72436
rect 11004 72382 11006 72434
rect 11006 72382 11058 72434
rect 11058 72382 11060 72434
rect 11004 72380 11060 72382
rect 10668 72044 10724 72100
rect 11116 72268 11172 72324
rect 10892 72044 10948 72100
rect 10668 71762 10724 71764
rect 10668 71710 10670 71762
rect 10670 71710 10722 71762
rect 10722 71710 10724 71762
rect 10668 71708 10724 71710
rect 10780 71260 10836 71316
rect 10892 71036 10948 71092
rect 10668 69692 10724 69748
rect 10444 68626 10500 68628
rect 10444 68574 10446 68626
rect 10446 68574 10498 68626
rect 10498 68574 10500 68626
rect 10444 68572 10500 68574
rect 10332 68348 10388 68404
rect 10332 68124 10388 68180
rect 10892 69186 10948 69188
rect 10892 69134 10894 69186
rect 10894 69134 10946 69186
rect 10946 69134 10948 69186
rect 10892 69132 10948 69134
rect 10780 68908 10836 68964
rect 11004 68796 11060 68852
rect 11116 70700 11172 70756
rect 10668 68572 10724 68628
rect 10892 68572 10948 68628
rect 10556 67228 10612 67284
rect 10668 67116 10724 67172
rect 10108 66892 10164 66948
rect 10556 66892 10612 66948
rect 10556 66274 10612 66276
rect 10556 66222 10558 66274
rect 10558 66222 10610 66274
rect 10610 66222 10612 66274
rect 10556 66220 10612 66222
rect 10444 65548 10500 65604
rect 10556 65884 10612 65940
rect 10220 65324 10276 65380
rect 10108 64988 10164 65044
rect 10108 64540 10164 64596
rect 9548 63644 9604 63700
rect 9996 63922 10052 63924
rect 9996 63870 9998 63922
rect 9998 63870 10050 63922
rect 10050 63870 10052 63922
rect 9996 63868 10052 63870
rect 9212 63138 9268 63140
rect 9212 63086 9214 63138
rect 9214 63086 9266 63138
rect 9266 63086 9268 63138
rect 9212 63084 9268 63086
rect 9324 62914 9380 62916
rect 9324 62862 9326 62914
rect 9326 62862 9378 62914
rect 9378 62862 9380 62914
rect 9324 62860 9380 62862
rect 9100 60172 9156 60228
rect 9212 62188 9268 62244
rect 8988 60114 9044 60116
rect 8988 60062 8990 60114
rect 8990 60062 9042 60114
rect 9042 60062 9044 60114
rect 8988 60060 9044 60062
rect 8652 59500 8708 59556
rect 9100 59442 9156 59444
rect 9100 59390 9102 59442
rect 9102 59390 9154 59442
rect 9154 59390 9156 59442
rect 9100 59388 9156 59390
rect 8988 59276 9044 59332
rect 9548 61964 9604 62020
rect 9436 60114 9492 60116
rect 9436 60062 9438 60114
rect 9438 60062 9490 60114
rect 9490 60062 9492 60114
rect 9436 60060 9492 60062
rect 9996 63420 10052 63476
rect 10332 65212 10388 65268
rect 10332 64988 10388 65044
rect 10444 64764 10500 64820
rect 10332 63810 10388 63812
rect 10332 63758 10334 63810
rect 10334 63758 10386 63810
rect 10386 63758 10388 63810
rect 10332 63756 10388 63758
rect 9996 63250 10052 63252
rect 9996 63198 9998 63250
rect 9998 63198 10050 63250
rect 10050 63198 10052 63250
rect 9996 63196 10052 63198
rect 10108 63084 10164 63140
rect 11004 68402 11060 68404
rect 11004 68350 11006 68402
rect 11006 68350 11058 68402
rect 11058 68350 11060 68402
rect 11004 68348 11060 68350
rect 10780 63084 10836 63140
rect 11452 74284 11508 74340
rect 11340 73948 11396 74004
rect 11340 73612 11396 73668
rect 11340 72492 11396 72548
rect 11452 73276 11508 73332
rect 10892 66444 10948 66500
rect 11340 71708 11396 71764
rect 11788 74396 11844 74452
rect 11788 73948 11844 74004
rect 12124 76636 12180 76692
rect 12124 75852 12180 75908
rect 12236 77420 12292 77476
rect 13804 77308 13860 77364
rect 12348 75852 12404 75908
rect 13580 76300 13636 76356
rect 13468 75852 13524 75908
rect 12908 75794 12964 75796
rect 12908 75742 12910 75794
rect 12910 75742 12962 75794
rect 12962 75742 12964 75794
rect 12908 75740 12964 75742
rect 13132 75068 13188 75124
rect 13020 75010 13076 75012
rect 13020 74958 13022 75010
rect 13022 74958 13074 75010
rect 13074 74958 13076 75010
rect 13020 74956 13076 74958
rect 12460 74620 12516 74676
rect 12012 74114 12068 74116
rect 12012 74062 12014 74114
rect 12014 74062 12066 74114
rect 12066 74062 12068 74114
rect 12012 74060 12068 74062
rect 11900 73836 11956 73892
rect 11788 73218 11844 73220
rect 11788 73166 11790 73218
rect 11790 73166 11842 73218
rect 11842 73166 11844 73218
rect 11788 73164 11844 73166
rect 11676 72828 11732 72884
rect 11564 72268 11620 72324
rect 11452 70252 11508 70308
rect 11676 71596 11732 71652
rect 11228 67730 11284 67732
rect 11228 67678 11230 67730
rect 11230 67678 11282 67730
rect 11282 67678 11284 67730
rect 11228 67676 11284 67678
rect 11900 72940 11956 72996
rect 12124 73948 12180 74004
rect 11900 71820 11956 71876
rect 11788 70700 11844 70756
rect 11676 69298 11732 69300
rect 11676 69246 11678 69298
rect 11678 69246 11730 69298
rect 11730 69246 11732 69298
rect 11676 69244 11732 69246
rect 11564 68796 11620 68852
rect 11340 66892 11396 66948
rect 11452 68236 11508 68292
rect 11676 68236 11732 68292
rect 11900 68236 11956 68292
rect 11788 67730 11844 67732
rect 11788 67678 11790 67730
rect 11790 67678 11842 67730
rect 11842 67678 11844 67730
rect 11788 67676 11844 67678
rect 11452 66668 11508 66724
rect 11116 66332 11172 66388
rect 11564 66162 11620 66164
rect 11564 66110 11566 66162
rect 11566 66110 11618 66162
rect 11618 66110 11620 66162
rect 11564 66108 11620 66110
rect 11228 65490 11284 65492
rect 11228 65438 11230 65490
rect 11230 65438 11282 65490
rect 11282 65438 11284 65490
rect 11228 65436 11284 65438
rect 10556 62972 10612 63028
rect 10220 62636 10276 62692
rect 10780 62578 10836 62580
rect 10780 62526 10782 62578
rect 10782 62526 10834 62578
rect 10834 62526 10836 62578
rect 10780 62524 10836 62526
rect 10668 62412 10724 62468
rect 9996 62242 10052 62244
rect 9996 62190 9998 62242
rect 9998 62190 10050 62242
rect 10050 62190 10052 62242
rect 9996 62188 10052 62190
rect 9772 62076 9828 62132
rect 10668 62242 10724 62244
rect 10668 62190 10670 62242
rect 10670 62190 10722 62242
rect 10722 62190 10724 62242
rect 10668 62188 10724 62190
rect 11452 64204 11508 64260
rect 11228 63868 11284 63924
rect 11340 63756 11396 63812
rect 11340 63308 11396 63364
rect 11564 63308 11620 63364
rect 11900 65324 11956 65380
rect 12236 72546 12292 72548
rect 12236 72494 12238 72546
rect 12238 72494 12290 72546
rect 12290 72494 12292 72546
rect 12236 72492 12292 72494
rect 13356 74786 13412 74788
rect 13356 74734 13358 74786
rect 13358 74734 13410 74786
rect 13410 74734 13412 74786
rect 13356 74732 13412 74734
rect 13132 74620 13188 74676
rect 12796 74002 12852 74004
rect 12796 73950 12798 74002
rect 12798 73950 12850 74002
rect 12850 73950 12852 74002
rect 12796 73948 12852 73950
rect 12796 73218 12852 73220
rect 12796 73166 12798 73218
rect 12798 73166 12850 73218
rect 12850 73166 12852 73218
rect 12796 73164 12852 73166
rect 12572 73052 12628 73108
rect 13020 73330 13076 73332
rect 13020 73278 13022 73330
rect 13022 73278 13074 73330
rect 13074 73278 13076 73330
rect 13020 73276 13076 73278
rect 12908 72380 12964 72436
rect 12684 71260 12740 71316
rect 12572 70924 12628 70980
rect 12460 70588 12516 70644
rect 13020 70924 13076 70980
rect 12908 70754 12964 70756
rect 12908 70702 12910 70754
rect 12910 70702 12962 70754
rect 12962 70702 12964 70754
rect 12908 70700 12964 70702
rect 12684 70588 12740 70644
rect 12124 69468 12180 69524
rect 12124 69132 12180 69188
rect 12684 69468 12740 69524
rect 12572 69020 12628 69076
rect 12236 66946 12292 66948
rect 12236 66894 12238 66946
rect 12238 66894 12290 66946
rect 12290 66894 12292 66946
rect 12236 66892 12292 66894
rect 12124 64652 12180 64708
rect 12684 68572 12740 68628
rect 12908 68572 12964 68628
rect 12684 67900 12740 67956
rect 12572 67340 12628 67396
rect 12684 67004 12740 67060
rect 12796 67228 12852 67284
rect 12796 66050 12852 66052
rect 12796 65998 12798 66050
rect 12798 65998 12850 66050
rect 12850 65998 12852 66050
rect 12796 65996 12852 65998
rect 12460 65660 12516 65716
rect 12348 64540 12404 64596
rect 12572 64428 12628 64484
rect 11900 63868 11956 63924
rect 11116 62748 11172 62804
rect 11788 63532 11844 63588
rect 11228 62354 11284 62356
rect 11228 62302 11230 62354
rect 11230 62302 11282 62354
rect 11282 62302 11284 62354
rect 11228 62300 11284 62302
rect 10556 61852 10612 61908
rect 10780 62076 10836 62132
rect 9884 61682 9940 61684
rect 9884 61630 9886 61682
rect 9886 61630 9938 61682
rect 9938 61630 9940 61682
rect 9884 61628 9940 61630
rect 10780 61682 10836 61684
rect 10780 61630 10782 61682
rect 10782 61630 10834 61682
rect 10834 61630 10836 61682
rect 10780 61628 10836 61630
rect 10220 61570 10276 61572
rect 10220 61518 10222 61570
rect 10222 61518 10274 61570
rect 10274 61518 10276 61570
rect 10220 61516 10276 61518
rect 11116 61570 11172 61572
rect 11116 61518 11118 61570
rect 11118 61518 11170 61570
rect 11170 61518 11172 61570
rect 11116 61516 11172 61518
rect 9772 60732 9828 60788
rect 9884 61404 9940 61460
rect 10108 61068 10164 61124
rect 10220 61010 10276 61012
rect 10220 60958 10222 61010
rect 10222 60958 10274 61010
rect 10274 60958 10276 61010
rect 10220 60956 10276 60958
rect 10780 61010 10836 61012
rect 10780 60958 10782 61010
rect 10782 60958 10834 61010
rect 10834 60958 10836 61010
rect 10780 60956 10836 60958
rect 11116 60956 11172 61012
rect 9884 60508 9940 60564
rect 10668 60508 10724 60564
rect 9996 59890 10052 59892
rect 9996 59838 9998 59890
rect 9998 59838 10050 59890
rect 10050 59838 10052 59890
rect 9996 59836 10052 59838
rect 9772 59164 9828 59220
rect 9324 58716 9380 58772
rect 8988 57874 9044 57876
rect 8988 57822 8990 57874
rect 8990 57822 9042 57874
rect 9042 57822 9044 57874
rect 8988 57820 9044 57822
rect 10556 59612 10612 59668
rect 10444 59164 10500 59220
rect 10220 59052 10276 59108
rect 8764 57708 8820 57764
rect 10220 57484 10276 57540
rect 8204 57036 8260 57092
rect 9996 57036 10052 57092
rect 9324 56978 9380 56980
rect 9324 56926 9326 56978
rect 9326 56926 9378 56978
rect 9378 56926 9380 56978
rect 9324 56924 9380 56926
rect 9772 56978 9828 56980
rect 9772 56926 9774 56978
rect 9774 56926 9826 56978
rect 9826 56926 9828 56978
rect 9772 56924 9828 56926
rect 9324 56700 9380 56756
rect 8092 55244 8148 55300
rect 7756 53676 7812 53732
rect 8316 53676 8372 53732
rect 7420 45164 7476 45220
rect 8204 45164 8260 45220
rect 5964 43596 6020 43652
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4284 41804 4340 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 8316 5964 8372 6020
rect 10780 59106 10836 59108
rect 10780 59054 10782 59106
rect 10782 59054 10834 59106
rect 10834 59054 10836 59106
rect 10780 59052 10836 59054
rect 10668 58434 10724 58436
rect 10668 58382 10670 58434
rect 10670 58382 10722 58434
rect 10722 58382 10724 58434
rect 10668 58380 10724 58382
rect 11228 60172 11284 60228
rect 11228 59442 11284 59444
rect 11228 59390 11230 59442
rect 11230 59390 11282 59442
rect 11282 59390 11284 59442
rect 11228 59388 11284 59390
rect 11564 62748 11620 62804
rect 12348 63756 12404 63812
rect 12012 63532 12068 63588
rect 12236 63138 12292 63140
rect 12236 63086 12238 63138
rect 12238 63086 12290 63138
rect 12290 63086 12292 63138
rect 12236 63084 12292 63086
rect 11900 62636 11956 62692
rect 12012 61516 12068 61572
rect 12124 62860 12180 62916
rect 11900 61404 11956 61460
rect 11340 59052 11396 59108
rect 11452 60396 11508 60452
rect 11452 59388 11508 59444
rect 11452 58940 11508 58996
rect 11900 60508 11956 60564
rect 12012 61346 12068 61348
rect 12012 61294 12014 61346
rect 12014 61294 12066 61346
rect 12066 61294 12068 61346
rect 12012 61292 12068 61294
rect 11564 60060 11620 60116
rect 11676 60172 11732 60228
rect 12572 63922 12628 63924
rect 12572 63870 12574 63922
rect 12574 63870 12626 63922
rect 12626 63870 12628 63922
rect 12572 63868 12628 63870
rect 12348 61516 12404 61572
rect 12908 67004 12964 67060
rect 13020 65436 13076 65492
rect 13356 74172 13412 74228
rect 13244 72268 13300 72324
rect 13804 75964 13860 76020
rect 13916 75852 13972 75908
rect 13692 75516 13748 75572
rect 14028 75628 14084 75684
rect 13804 75458 13860 75460
rect 13804 75406 13806 75458
rect 13806 75406 13858 75458
rect 13858 75406 13860 75458
rect 13804 75404 13860 75406
rect 13692 75292 13748 75348
rect 13468 71708 13524 71764
rect 14140 74060 14196 74116
rect 13244 71148 13300 71204
rect 13356 71650 13412 71652
rect 13356 71598 13358 71650
rect 13358 71598 13410 71650
rect 13410 71598 13412 71650
rect 13356 71596 13412 71598
rect 13468 71484 13524 71540
rect 13692 71484 13748 71540
rect 13804 71932 13860 71988
rect 13580 71260 13636 71316
rect 14028 71596 14084 71652
rect 14252 72716 14308 72772
rect 14476 79660 14532 79716
rect 15148 79324 15204 79380
rect 14588 77868 14644 77924
rect 14364 73836 14420 73892
rect 13916 71260 13972 71316
rect 14028 71148 14084 71204
rect 14476 71820 14532 71876
rect 13804 71036 13860 71092
rect 13692 70700 13748 70756
rect 13468 69692 13524 69748
rect 13468 68908 13524 68964
rect 12908 64652 12964 64708
rect 12908 63980 12964 64036
rect 12796 62860 12852 62916
rect 13020 62636 13076 62692
rect 13132 64092 13188 64148
rect 12684 61740 12740 61796
rect 12908 61964 12964 62020
rect 12348 60508 12404 60564
rect 12124 60284 12180 60340
rect 12012 60172 12068 60228
rect 12684 60508 12740 60564
rect 12796 60060 12852 60116
rect 13020 60508 13076 60564
rect 12796 59612 12852 59668
rect 12908 59724 12964 59780
rect 12124 58546 12180 58548
rect 12124 58494 12126 58546
rect 12126 58494 12178 58546
rect 12178 58494 12180 58546
rect 12124 58492 12180 58494
rect 12572 58546 12628 58548
rect 12572 58494 12574 58546
rect 12574 58494 12626 58546
rect 12626 58494 12628 58546
rect 12572 58492 12628 58494
rect 12012 58156 12068 58212
rect 11564 57874 11620 57876
rect 11564 57822 11566 57874
rect 11566 57822 11618 57874
rect 11618 57822 11620 57874
rect 11564 57820 11620 57822
rect 12460 57874 12516 57876
rect 12460 57822 12462 57874
rect 12462 57822 12514 57874
rect 12514 57822 12516 57874
rect 12460 57820 12516 57822
rect 12460 57596 12516 57652
rect 10332 51996 10388 52052
rect 11676 56588 11732 56644
rect 11676 50316 11732 50372
rect 9996 48300 10052 48356
rect 8204 5852 8260 5908
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6972 3612 7028 3668
rect 3500 3554 3556 3556
rect 3500 3502 3502 3554
rect 3502 3502 3554 3554
rect 3554 3502 3556 3554
rect 3500 3500 3556 3502
rect 4284 3554 4340 3556
rect 4284 3502 4286 3554
rect 4286 3502 4338 3554
rect 4338 3502 4340 3554
rect 4284 3500 4340 3502
rect 11004 6076 11060 6132
rect 17948 79436 18004 79492
rect 15932 78764 15988 78820
rect 17388 78876 17444 78932
rect 15932 76188 15988 76244
rect 15148 74396 15204 74452
rect 14812 73500 14868 73556
rect 15036 72380 15092 72436
rect 14588 70700 14644 70756
rect 13692 70252 13748 70308
rect 13692 69356 13748 69412
rect 13804 67788 13860 67844
rect 13692 66386 13748 66388
rect 13692 66334 13694 66386
rect 13694 66334 13746 66386
rect 13746 66334 13748 66386
rect 13692 66332 13748 66334
rect 13804 65324 13860 65380
rect 13580 64876 13636 64932
rect 13468 64764 13524 64820
rect 13916 64652 13972 64708
rect 13916 64428 13972 64484
rect 13580 64204 13636 64260
rect 13356 62748 13412 62804
rect 13356 62412 13412 62468
rect 13692 64092 13748 64148
rect 14028 68066 14084 68068
rect 14028 68014 14030 68066
rect 14030 68014 14082 68066
rect 14082 68014 14084 68066
rect 14028 68012 14084 68014
rect 14028 64092 14084 64148
rect 14924 70588 14980 70644
rect 14812 67788 14868 67844
rect 14252 67004 14308 67060
rect 14476 67004 14532 67060
rect 14364 66946 14420 66948
rect 14364 66894 14366 66946
rect 14366 66894 14418 66946
rect 14418 66894 14420 66946
rect 14364 66892 14420 66894
rect 14588 66556 14644 66612
rect 14364 66108 14420 66164
rect 14252 64930 14308 64932
rect 14252 64878 14254 64930
rect 14254 64878 14306 64930
rect 14306 64878 14308 64930
rect 14252 64876 14308 64878
rect 15484 75964 15540 76020
rect 15372 71148 15428 71204
rect 15260 70812 15316 70868
rect 15148 68796 15204 68852
rect 15372 70588 15428 70644
rect 15148 67058 15204 67060
rect 15148 67006 15150 67058
rect 15150 67006 15202 67058
rect 15202 67006 15204 67058
rect 15148 67004 15204 67006
rect 16716 76466 16772 76468
rect 16716 76414 16718 76466
rect 16718 76414 16770 76466
rect 16770 76414 16772 76466
rect 16716 76412 16772 76414
rect 16828 75794 16884 75796
rect 16828 75742 16830 75794
rect 16830 75742 16882 75794
rect 16882 75742 16884 75794
rect 16828 75740 16884 75742
rect 16044 74956 16100 75012
rect 16940 75628 16996 75684
rect 17500 75682 17556 75684
rect 17500 75630 17502 75682
rect 17502 75630 17554 75682
rect 17554 75630 17556 75682
rect 17500 75628 17556 75630
rect 17724 75068 17780 75124
rect 16604 74284 16660 74340
rect 16716 72434 16772 72436
rect 16716 72382 16718 72434
rect 16718 72382 16770 72434
rect 16770 72382 16772 72434
rect 16716 72380 16772 72382
rect 16380 70588 16436 70644
rect 16716 70588 16772 70644
rect 16492 70476 16548 70532
rect 16156 69916 16212 69972
rect 15596 68348 15652 68404
rect 15708 67954 15764 67956
rect 15708 67902 15710 67954
rect 15710 67902 15762 67954
rect 15762 67902 15764 67954
rect 15708 67900 15764 67902
rect 15596 67340 15652 67396
rect 15596 67058 15652 67060
rect 15596 67006 15598 67058
rect 15598 67006 15650 67058
rect 15650 67006 15652 67058
rect 15596 67004 15652 67006
rect 14812 66108 14868 66164
rect 15036 66332 15092 66388
rect 14812 65490 14868 65492
rect 14812 65438 14814 65490
rect 14814 65438 14866 65490
rect 14866 65438 14868 65490
rect 14812 65436 14868 65438
rect 15036 64652 15092 64708
rect 16604 69692 16660 69748
rect 16492 68908 16548 68964
rect 16380 68236 16436 68292
rect 16268 67842 16324 67844
rect 16268 67790 16270 67842
rect 16270 67790 16322 67842
rect 16322 67790 16324 67842
rect 16268 67788 16324 67790
rect 15820 67228 15876 67284
rect 15932 67564 15988 67620
rect 15708 66220 15764 66276
rect 15820 65772 15876 65828
rect 15596 65490 15652 65492
rect 15596 65438 15598 65490
rect 15598 65438 15650 65490
rect 15650 65438 15652 65490
rect 15596 65436 15652 65438
rect 15932 64988 15988 65044
rect 16044 65996 16100 66052
rect 15372 64930 15428 64932
rect 15372 64878 15374 64930
rect 15374 64878 15426 64930
rect 15426 64878 15428 64930
rect 15372 64876 15428 64878
rect 15260 64204 15316 64260
rect 13692 63026 13748 63028
rect 13692 62974 13694 63026
rect 13694 62974 13746 63026
rect 13746 62974 13748 63026
rect 13692 62972 13748 62974
rect 13692 62748 13748 62804
rect 13356 61740 13412 61796
rect 13580 62354 13636 62356
rect 13580 62302 13582 62354
rect 13582 62302 13634 62354
rect 13634 62302 13636 62354
rect 13580 62300 13636 62302
rect 13692 61964 13748 62020
rect 13804 61852 13860 61908
rect 14364 63138 14420 63140
rect 14364 63086 14366 63138
rect 14366 63086 14418 63138
rect 14418 63086 14420 63138
rect 14364 63084 14420 63086
rect 14028 62188 14084 62244
rect 14364 62076 14420 62132
rect 13916 61628 13972 61684
rect 14140 61852 14196 61908
rect 13692 61346 13748 61348
rect 13692 61294 13694 61346
rect 13694 61294 13746 61346
rect 13746 61294 13748 61346
rect 13692 61292 13748 61294
rect 13916 61180 13972 61236
rect 13692 61010 13748 61012
rect 13692 60958 13694 61010
rect 13694 60958 13746 61010
rect 13746 60958 13748 61010
rect 13692 60956 13748 60958
rect 13468 60844 13524 60900
rect 14028 60898 14084 60900
rect 14028 60846 14030 60898
rect 14030 60846 14082 60898
rect 14082 60846 14084 60898
rect 14028 60844 14084 60846
rect 13916 60508 13972 60564
rect 14364 61852 14420 61908
rect 14700 61458 14756 61460
rect 14700 61406 14702 61458
rect 14702 61406 14754 61458
rect 14754 61406 14756 61458
rect 14700 61404 14756 61406
rect 14252 61068 14308 61124
rect 14364 61292 14420 61348
rect 14140 60172 14196 60228
rect 13356 60060 13412 60116
rect 13580 59330 13636 59332
rect 13580 59278 13582 59330
rect 13582 59278 13634 59330
rect 13634 59278 13636 59330
rect 13580 59276 13636 59278
rect 13692 58546 13748 58548
rect 13692 58494 13694 58546
rect 13694 58494 13746 58546
rect 13746 58494 13748 58546
rect 13692 58492 13748 58494
rect 13804 57762 13860 57764
rect 13804 57710 13806 57762
rect 13806 57710 13858 57762
rect 13858 57710 13860 57762
rect 13804 57708 13860 57710
rect 13356 57538 13412 57540
rect 13356 57486 13358 57538
rect 13358 57486 13410 57538
rect 13410 57486 13412 57538
rect 13356 57484 13412 57486
rect 13580 56866 13636 56868
rect 13580 56814 13582 56866
rect 13582 56814 13634 56866
rect 13634 56814 13636 56866
rect 13580 56812 13636 56814
rect 12908 56642 12964 56644
rect 12908 56590 12910 56642
rect 12910 56590 12962 56642
rect 12962 56590 12964 56642
rect 12908 56588 12964 56590
rect 12572 56476 12628 56532
rect 14028 57484 14084 57540
rect 14252 60844 14308 60900
rect 15148 64146 15204 64148
rect 15148 64094 15150 64146
rect 15150 64094 15202 64146
rect 15202 64094 15204 64146
rect 15148 64092 15204 64094
rect 15484 63922 15540 63924
rect 15484 63870 15486 63922
rect 15486 63870 15538 63922
rect 15538 63870 15540 63922
rect 15484 63868 15540 63870
rect 15260 63420 15316 63476
rect 15260 63250 15316 63252
rect 15260 63198 15262 63250
rect 15262 63198 15314 63250
rect 15314 63198 15316 63250
rect 15260 63196 15316 63198
rect 15708 63980 15764 64036
rect 15932 64706 15988 64708
rect 15932 64654 15934 64706
rect 15934 64654 15986 64706
rect 15986 64654 15988 64706
rect 15932 64652 15988 64654
rect 16044 64428 16100 64484
rect 16044 63420 16100 63476
rect 15708 63196 15764 63252
rect 15596 63084 15652 63140
rect 15260 62972 15316 63028
rect 15596 62636 15652 62692
rect 15260 62578 15316 62580
rect 15260 62526 15262 62578
rect 15262 62526 15314 62578
rect 15314 62526 15316 62578
rect 15260 62524 15316 62526
rect 14924 61404 14980 61460
rect 15036 61628 15092 61684
rect 15148 61570 15204 61572
rect 15148 61518 15150 61570
rect 15150 61518 15202 61570
rect 15202 61518 15204 61570
rect 15148 61516 15204 61518
rect 14924 60844 14980 60900
rect 15036 60732 15092 60788
rect 15372 59890 15428 59892
rect 15372 59838 15374 59890
rect 15374 59838 15426 59890
rect 15426 59838 15428 59890
rect 15372 59836 15428 59838
rect 15484 59442 15540 59444
rect 15484 59390 15486 59442
rect 15486 59390 15538 59442
rect 15538 59390 15540 59442
rect 15484 59388 15540 59390
rect 15820 62636 15876 62692
rect 15708 62130 15764 62132
rect 15708 62078 15710 62130
rect 15710 62078 15762 62130
rect 15762 62078 15764 62130
rect 15708 62076 15764 62078
rect 16044 62076 16100 62132
rect 15932 61964 15988 62020
rect 15708 61794 15764 61796
rect 15708 61742 15710 61794
rect 15710 61742 15762 61794
rect 15762 61742 15764 61794
rect 15708 61740 15764 61742
rect 15372 58546 15428 58548
rect 15372 58494 15374 58546
rect 15374 58494 15426 58546
rect 15426 58494 15428 58546
rect 15372 58492 15428 58494
rect 14476 58210 14532 58212
rect 14476 58158 14478 58210
rect 14478 58158 14530 58210
rect 14530 58158 14532 58210
rect 14476 58156 14532 58158
rect 14252 57650 14308 57652
rect 14252 57598 14254 57650
rect 14254 57598 14306 57650
rect 14306 57598 14308 57650
rect 14252 57596 14308 57598
rect 14700 57820 14756 57876
rect 15148 57874 15204 57876
rect 15148 57822 15150 57874
rect 15150 57822 15202 57874
rect 15202 57822 15204 57874
rect 15148 57820 15204 57822
rect 14700 57538 14756 57540
rect 14700 57486 14702 57538
rect 14702 57486 14754 57538
rect 14754 57486 14756 57538
rect 14700 57484 14756 57486
rect 14476 56252 14532 56308
rect 15148 56812 15204 56868
rect 16604 69132 16660 69188
rect 16940 70476 16996 70532
rect 16716 67676 16772 67732
rect 16604 67058 16660 67060
rect 16604 67006 16606 67058
rect 16606 67006 16658 67058
rect 16658 67006 16660 67058
rect 16604 67004 16660 67006
rect 16604 66668 16660 66724
rect 16828 67228 16884 67284
rect 17500 74732 17556 74788
rect 17164 69692 17220 69748
rect 17388 71820 17444 71876
rect 17388 70028 17444 70084
rect 16940 67116 16996 67172
rect 16940 66946 16996 66948
rect 16940 66894 16942 66946
rect 16942 66894 16994 66946
rect 16994 66894 16996 66946
rect 16940 66892 16996 66894
rect 16268 65602 16324 65604
rect 16268 65550 16270 65602
rect 16270 65550 16322 65602
rect 16322 65550 16324 65602
rect 16268 65548 16324 65550
rect 16604 65490 16660 65492
rect 16604 65438 16606 65490
rect 16606 65438 16658 65490
rect 16658 65438 16660 65490
rect 16604 65436 16660 65438
rect 16268 65378 16324 65380
rect 16268 65326 16270 65378
rect 16270 65326 16322 65378
rect 16322 65326 16324 65378
rect 16268 65324 16324 65326
rect 16716 65212 16772 65268
rect 16380 64540 16436 64596
rect 16492 64988 16548 65044
rect 16604 64428 16660 64484
rect 17164 67954 17220 67956
rect 17164 67902 17166 67954
rect 17166 67902 17218 67954
rect 17218 67902 17220 67954
rect 17164 67900 17220 67902
rect 17724 73330 17780 73332
rect 17724 73278 17726 73330
rect 17726 73278 17778 73330
rect 17778 73278 17780 73330
rect 17724 73276 17780 73278
rect 28812 79660 28868 79716
rect 28364 79548 28420 79604
rect 18396 79100 18452 79156
rect 18060 76076 18116 76132
rect 18732 78988 18788 79044
rect 18508 76354 18564 76356
rect 18508 76302 18510 76354
rect 18510 76302 18562 76354
rect 18562 76302 18564 76354
rect 18508 76300 18564 76302
rect 18620 75852 18676 75908
rect 18172 75292 18228 75348
rect 17724 73052 17780 73108
rect 17612 70700 17668 70756
rect 18396 75458 18452 75460
rect 18396 75406 18398 75458
rect 18398 75406 18450 75458
rect 18450 75406 18452 75458
rect 18396 75404 18452 75406
rect 18396 74508 18452 74564
rect 20412 78540 20468 78596
rect 20188 78092 20244 78148
rect 19068 77980 19124 78036
rect 18844 76524 18900 76580
rect 18732 75010 18788 75012
rect 18732 74958 18734 75010
rect 18734 74958 18786 75010
rect 18786 74958 18788 75010
rect 18732 74956 18788 74958
rect 18620 74508 18676 74564
rect 18508 73442 18564 73444
rect 18508 73390 18510 73442
rect 18510 73390 18562 73442
rect 18562 73390 18564 73442
rect 18508 73388 18564 73390
rect 18396 73106 18452 73108
rect 18396 73054 18398 73106
rect 18398 73054 18450 73106
rect 18450 73054 18452 73106
rect 18396 73052 18452 73054
rect 18396 72492 18452 72548
rect 18172 72380 18228 72436
rect 18060 71986 18116 71988
rect 18060 71934 18062 71986
rect 18062 71934 18114 71986
rect 18114 71934 18116 71986
rect 18060 71932 18116 71934
rect 17948 69804 18004 69860
rect 18396 70924 18452 70980
rect 18508 72268 18564 72324
rect 18396 70140 18452 70196
rect 18396 69916 18452 69972
rect 18172 69580 18228 69636
rect 18284 69804 18340 69860
rect 18060 69020 18116 69076
rect 17836 68684 17892 68740
rect 18172 68684 18228 68740
rect 18508 69580 18564 69636
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19404 75516 19460 75572
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 20300 76412 20356 76468
rect 20300 75628 20356 75684
rect 18956 72940 19012 72996
rect 18732 71596 18788 71652
rect 18844 70476 18900 70532
rect 18620 69356 18676 69412
rect 18508 68236 18564 68292
rect 17836 68012 17892 68068
rect 17724 67564 17780 67620
rect 18620 67788 18676 67844
rect 17500 67228 17556 67284
rect 17948 67282 18004 67284
rect 17948 67230 17950 67282
rect 17950 67230 18002 67282
rect 18002 67230 18004 67282
rect 17948 67228 18004 67230
rect 17388 66892 17444 66948
rect 18284 67058 18340 67060
rect 18284 67006 18286 67058
rect 18286 67006 18338 67058
rect 18338 67006 18340 67058
rect 18284 67004 18340 67006
rect 18732 67228 18788 67284
rect 18844 70028 18900 70084
rect 17836 66946 17892 66948
rect 17836 66894 17838 66946
rect 17838 66894 17890 66946
rect 17890 66894 17892 66946
rect 17836 66892 17892 66894
rect 17164 66556 17220 66612
rect 17164 64706 17220 64708
rect 17164 64654 17166 64706
rect 17166 64654 17218 64706
rect 17218 64654 17220 64706
rect 17164 64652 17220 64654
rect 17164 64428 17220 64484
rect 16604 63644 16660 63700
rect 16380 63196 16436 63252
rect 16828 64092 16884 64148
rect 17052 63980 17108 64036
rect 16716 63308 16772 63364
rect 16716 62972 16772 63028
rect 16716 62578 16772 62580
rect 16716 62526 16718 62578
rect 16718 62526 16770 62578
rect 16770 62526 16772 62578
rect 16716 62524 16772 62526
rect 16380 61964 16436 62020
rect 15820 61570 15876 61572
rect 15820 61518 15822 61570
rect 15822 61518 15874 61570
rect 15874 61518 15876 61570
rect 15820 61516 15876 61518
rect 16044 61404 16100 61460
rect 15820 60898 15876 60900
rect 15820 60846 15822 60898
rect 15822 60846 15874 60898
rect 15874 60846 15876 60898
rect 15820 60844 15876 60846
rect 16268 60172 16324 60228
rect 15820 60114 15876 60116
rect 15820 60062 15822 60114
rect 15822 60062 15874 60114
rect 15874 60062 15876 60114
rect 15820 60060 15876 60062
rect 16380 60284 16436 60340
rect 15932 59612 15988 59668
rect 15932 58716 15988 58772
rect 15708 55020 15764 55076
rect 16828 61964 16884 62020
rect 16716 61458 16772 61460
rect 16716 61406 16718 61458
rect 16718 61406 16770 61458
rect 16770 61406 16772 61458
rect 16716 61404 16772 61406
rect 16940 61628 16996 61684
rect 16940 61292 16996 61348
rect 17052 63756 17108 63812
rect 16828 60956 16884 61012
rect 17164 62412 17220 62468
rect 17164 62076 17220 62132
rect 18060 66556 18116 66612
rect 18284 66780 18340 66836
rect 18620 66220 18676 66276
rect 17836 66108 17892 66164
rect 17500 64876 17556 64932
rect 17948 66050 18004 66052
rect 17948 65998 17950 66050
rect 17950 65998 18002 66050
rect 18002 65998 18004 66050
rect 17948 65996 18004 65998
rect 18844 66668 18900 66724
rect 18732 66444 18788 66500
rect 17948 65660 18004 65716
rect 18172 65714 18228 65716
rect 18172 65662 18174 65714
rect 18174 65662 18226 65714
rect 18226 65662 18228 65714
rect 18172 65660 18228 65662
rect 17388 63644 17444 63700
rect 17612 64428 17668 64484
rect 17724 63810 17780 63812
rect 17724 63758 17726 63810
rect 17726 63758 17778 63810
rect 17778 63758 17780 63810
rect 17724 63756 17780 63758
rect 17612 62524 17668 62580
rect 17500 61964 17556 62020
rect 16828 60620 16884 60676
rect 17276 59778 17332 59780
rect 17276 59726 17278 59778
rect 17278 59726 17330 59778
rect 17330 59726 17332 59778
rect 17276 59724 17332 59726
rect 16940 59442 16996 59444
rect 16940 59390 16942 59442
rect 16942 59390 16994 59442
rect 16994 59390 16996 59442
rect 16940 59388 16996 59390
rect 16828 58940 16884 58996
rect 16716 58604 16772 58660
rect 16156 54908 16212 54964
rect 15148 41804 15204 41860
rect 15148 40348 15204 40404
rect 15932 40348 15988 40404
rect 13804 36652 13860 36708
rect 14812 6748 14868 6804
rect 12460 6130 12516 6132
rect 12460 6078 12462 6130
rect 12462 6078 12514 6130
rect 12514 6078 12516 6130
rect 12460 6076 12516 6078
rect 15036 5964 15092 6020
rect 11228 4508 11284 4564
rect 9996 4396 10052 4452
rect 7644 4338 7700 4340
rect 7644 4286 7646 4338
rect 7646 4286 7698 4338
rect 7698 4286 7700 4338
rect 7644 4284 7700 4286
rect 11340 4338 11396 4340
rect 11340 4286 11342 4338
rect 11342 4286 11394 4338
rect 11394 4286 11396 4338
rect 11340 4284 11396 4286
rect 7868 3666 7924 3668
rect 7868 3614 7870 3666
rect 7870 3614 7922 3666
rect 7922 3614 7924 3666
rect 7868 3612 7924 3614
rect 11676 4508 11732 4564
rect 12348 4562 12404 4564
rect 12348 4510 12350 4562
rect 12350 4510 12402 4562
rect 12402 4510 12404 4562
rect 12348 4508 12404 4510
rect 14588 4562 14644 4564
rect 14588 4510 14590 4562
rect 14590 4510 14642 4562
rect 14642 4510 14644 4562
rect 14588 4508 14644 4510
rect 11900 4396 11956 4452
rect 12796 4450 12852 4452
rect 12796 4398 12798 4450
rect 12798 4398 12850 4450
rect 12850 4398 12852 4450
rect 12796 4396 12852 4398
rect 15932 5964 15988 6020
rect 15372 5794 15428 5796
rect 15372 5742 15374 5794
rect 15374 5742 15426 5794
rect 15426 5742 15428 5794
rect 15372 5740 15428 5742
rect 17164 58604 17220 58660
rect 17612 60898 17668 60900
rect 17612 60846 17614 60898
rect 17614 60846 17666 60898
rect 17666 60846 17668 60898
rect 17612 60844 17668 60846
rect 18284 64764 18340 64820
rect 18508 64652 18564 64708
rect 18396 64594 18452 64596
rect 18396 64542 18398 64594
rect 18398 64542 18450 64594
rect 18450 64542 18452 64594
rect 18396 64540 18452 64542
rect 18172 64316 18228 64372
rect 18284 64092 18340 64148
rect 17948 62636 18004 62692
rect 18172 63868 18228 63924
rect 18396 63922 18452 63924
rect 18396 63870 18398 63922
rect 18398 63870 18450 63922
rect 18450 63870 18452 63922
rect 18396 63868 18452 63870
rect 18620 63644 18676 63700
rect 18732 64316 18788 64372
rect 18620 63308 18676 63364
rect 18060 61516 18116 61572
rect 18172 62300 18228 62356
rect 19180 70588 19236 70644
rect 24556 78428 24612 78484
rect 22988 78316 23044 78372
rect 20636 76524 20692 76580
rect 22316 76412 22372 76468
rect 21420 76354 21476 76356
rect 21420 76302 21422 76354
rect 21422 76302 21474 76354
rect 21474 76302 21476 76354
rect 21420 76300 21476 76302
rect 20076 74226 20132 74228
rect 20076 74174 20078 74226
rect 20078 74174 20130 74226
rect 20130 74174 20132 74226
rect 20076 74172 20132 74174
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19740 72940 19796 72996
rect 20300 72828 20356 72884
rect 19516 72322 19572 72324
rect 19516 72270 19518 72322
rect 19518 72270 19570 72322
rect 19570 72270 19572 72322
rect 19516 72268 19572 72270
rect 19404 72156 19460 72212
rect 19404 70924 19460 70980
rect 19516 70082 19572 70084
rect 19516 70030 19518 70082
rect 19518 70030 19570 70082
rect 19570 70030 19572 70082
rect 19516 70028 19572 70030
rect 23548 77308 23604 77364
rect 24332 76466 24388 76468
rect 24332 76414 24334 76466
rect 24334 76414 24386 76466
rect 24386 76414 24388 76466
rect 24332 76412 24388 76414
rect 22316 75682 22372 75684
rect 22316 75630 22318 75682
rect 22318 75630 22370 75682
rect 22370 75630 22372 75682
rect 22316 75628 22372 75630
rect 21756 74620 21812 74676
rect 21532 74060 21588 74116
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 20412 72268 20468 72324
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19628 69804 19684 69860
rect 20412 70364 20468 70420
rect 20188 70082 20244 70084
rect 20188 70030 20190 70082
rect 20190 70030 20242 70082
rect 20242 70030 20244 70082
rect 20188 70028 20244 70030
rect 19964 69132 20020 69188
rect 19836 69018 19892 69020
rect 19292 68908 19348 68964
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 20636 72434 20692 72436
rect 20636 72382 20638 72434
rect 20638 72382 20690 72434
rect 20690 72382 20692 72434
rect 20636 72380 20692 72382
rect 20188 68908 20244 68964
rect 20076 68124 20132 68180
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 20076 67170 20132 67172
rect 20076 67118 20078 67170
rect 20078 67118 20130 67170
rect 20130 67118 20132 67170
rect 20076 67116 20132 67118
rect 19964 66444 20020 66500
rect 19292 66386 19348 66388
rect 19292 66334 19294 66386
rect 19294 66334 19346 66386
rect 19346 66334 19348 66386
rect 19292 66332 19348 66334
rect 19068 65436 19124 65492
rect 19180 66220 19236 66276
rect 20076 66386 20132 66388
rect 20076 66334 20078 66386
rect 20078 66334 20130 66386
rect 20130 66334 20132 66386
rect 20076 66332 20132 66334
rect 20860 73218 20916 73220
rect 20860 73166 20862 73218
rect 20862 73166 20914 73218
rect 20914 73166 20916 73218
rect 20860 73164 20916 73166
rect 20860 71148 20916 71204
rect 20972 70700 21028 70756
rect 21084 73164 21140 73220
rect 21644 74002 21700 74004
rect 21644 73950 21646 74002
rect 21646 73950 21698 74002
rect 21698 73950 21700 74002
rect 21644 73948 21700 73950
rect 22092 74732 22148 74788
rect 21868 73890 21924 73892
rect 21868 73838 21870 73890
rect 21870 73838 21922 73890
rect 21922 73838 21924 73890
rect 21868 73836 21924 73838
rect 21756 72156 21812 72212
rect 20300 66220 20356 66276
rect 21644 70588 21700 70644
rect 20300 65996 20356 66052
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 20188 65772 20244 65828
rect 19628 65660 19684 65716
rect 19180 65100 19236 65156
rect 18956 64092 19012 64148
rect 18844 63980 18900 64036
rect 19740 64764 19796 64820
rect 19852 64428 19908 64484
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 17836 60060 17892 60116
rect 18172 61292 18228 61348
rect 17724 59724 17780 59780
rect 17724 58716 17780 58772
rect 17500 58380 17556 58436
rect 16828 55244 16884 55300
rect 18284 61010 18340 61012
rect 18284 60958 18286 61010
rect 18286 60958 18338 61010
rect 18338 60958 18340 61010
rect 18284 60956 18340 60958
rect 18956 63644 19012 63700
rect 18844 62076 18900 62132
rect 18732 61964 18788 62020
rect 18844 61180 18900 61236
rect 18508 60060 18564 60116
rect 18284 60002 18340 60004
rect 18284 59950 18286 60002
rect 18286 59950 18338 60002
rect 18338 59950 18340 60002
rect 18284 59948 18340 59950
rect 18060 59164 18116 59220
rect 18172 58940 18228 58996
rect 19292 63922 19348 63924
rect 19292 63870 19294 63922
rect 19294 63870 19346 63922
rect 19346 63870 19348 63922
rect 19292 63868 19348 63870
rect 19180 63756 19236 63812
rect 19292 62242 19348 62244
rect 19292 62190 19294 62242
rect 19294 62190 19346 62242
rect 19346 62190 19348 62242
rect 19292 62188 19348 62190
rect 19180 61068 19236 61124
rect 19068 60956 19124 61012
rect 19740 64092 19796 64148
rect 20300 64146 20356 64148
rect 20300 64094 20302 64146
rect 20302 64094 20354 64146
rect 20354 64094 20356 64146
rect 20300 64092 20356 64094
rect 20188 64034 20244 64036
rect 20188 63982 20190 64034
rect 20190 63982 20242 64034
rect 20242 63982 20244 64034
rect 20188 63980 20244 63982
rect 20300 63868 20356 63924
rect 22764 74002 22820 74004
rect 22764 73950 22766 74002
rect 22766 73950 22818 74002
rect 22818 73950 22820 74002
rect 22764 73948 22820 73950
rect 21308 69804 21364 69860
rect 20524 69298 20580 69300
rect 20524 69246 20526 69298
rect 20526 69246 20578 69298
rect 20578 69246 20580 69298
rect 20524 69244 20580 69246
rect 20972 69244 21028 69300
rect 21308 69244 21364 69300
rect 20748 69020 20804 69076
rect 21196 69020 21252 69076
rect 21196 68124 21252 68180
rect 20860 67452 20916 67508
rect 20860 66892 20916 66948
rect 20636 65996 20692 66052
rect 20748 66556 20804 66612
rect 20524 65266 20580 65268
rect 20524 65214 20526 65266
rect 20526 65214 20578 65266
rect 20578 65214 20580 65266
rect 20524 65212 20580 65214
rect 20524 64818 20580 64820
rect 20524 64766 20526 64818
rect 20526 64766 20578 64818
rect 20578 64766 20580 64818
rect 20524 64764 20580 64766
rect 19516 62300 19572 62356
rect 19180 60396 19236 60452
rect 19068 59890 19124 59892
rect 19068 59838 19070 59890
rect 19070 59838 19122 59890
rect 19122 59838 19124 59890
rect 19068 59836 19124 59838
rect 18844 59276 18900 59332
rect 18956 58492 19012 58548
rect 19740 63026 19796 63028
rect 19740 62974 19742 63026
rect 19742 62974 19794 63026
rect 19794 62974 19796 63026
rect 19740 62972 19796 62974
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19740 62578 19796 62580
rect 19740 62526 19742 62578
rect 19742 62526 19794 62578
rect 19794 62526 19796 62578
rect 19740 62524 19796 62526
rect 20412 63250 20468 63252
rect 20412 63198 20414 63250
rect 20414 63198 20466 63250
rect 20466 63198 20468 63250
rect 20412 63196 20468 63198
rect 19628 62188 19684 62244
rect 19740 61570 19796 61572
rect 19740 61518 19742 61570
rect 19742 61518 19794 61570
rect 19794 61518 19796 61570
rect 19740 61516 19796 61518
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19740 61010 19796 61012
rect 19740 60958 19742 61010
rect 19742 60958 19794 61010
rect 19794 60958 19796 61010
rect 19740 60956 19796 60958
rect 20412 61852 20468 61908
rect 20300 61346 20356 61348
rect 20300 61294 20302 61346
rect 20302 61294 20354 61346
rect 20354 61294 20356 61346
rect 20300 61292 20356 61294
rect 20188 60674 20244 60676
rect 20188 60622 20190 60674
rect 20190 60622 20242 60674
rect 20242 60622 20244 60674
rect 20188 60620 20244 60622
rect 20636 63644 20692 63700
rect 20860 65660 20916 65716
rect 20972 65548 21028 65604
rect 20860 64092 20916 64148
rect 20860 62914 20916 62916
rect 20860 62862 20862 62914
rect 20862 62862 20914 62914
rect 20914 62862 20916 62914
rect 20860 62860 20916 62862
rect 20860 62636 20916 62692
rect 20860 62300 20916 62356
rect 21196 64540 21252 64596
rect 21756 68796 21812 68852
rect 22988 73218 23044 73220
rect 22988 73166 22990 73218
rect 22990 73166 23042 73218
rect 23042 73166 23044 73218
rect 22988 73164 23044 73166
rect 21868 68348 21924 68404
rect 22652 71260 22708 71316
rect 21308 63980 21364 64036
rect 21420 67788 21476 67844
rect 21756 67842 21812 67844
rect 21756 67790 21758 67842
rect 21758 67790 21810 67842
rect 21810 67790 21812 67842
rect 21756 67788 21812 67790
rect 21644 67340 21700 67396
rect 21532 67228 21588 67284
rect 21868 66444 21924 66500
rect 21756 65996 21812 66052
rect 21868 65884 21924 65940
rect 21868 65548 21924 65604
rect 22428 69468 22484 69524
rect 22540 69692 22596 69748
rect 22204 69132 22260 69188
rect 22092 67004 22148 67060
rect 21532 64876 21588 64932
rect 22092 66332 22148 66388
rect 21308 63644 21364 63700
rect 21532 62860 21588 62916
rect 21756 63196 21812 63252
rect 22092 64540 22148 64596
rect 21980 63308 22036 63364
rect 21868 63138 21924 63140
rect 21868 63086 21870 63138
rect 21870 63086 21922 63138
rect 21922 63086 21924 63138
rect 21868 63084 21924 63086
rect 22204 64092 22260 64148
rect 22876 70588 22932 70644
rect 22652 67004 22708 67060
rect 22764 70140 22820 70196
rect 22764 66556 22820 66612
rect 22540 65884 22596 65940
rect 22652 66332 22708 66388
rect 22540 65602 22596 65604
rect 22540 65550 22542 65602
rect 22542 65550 22594 65602
rect 22594 65550 22596 65602
rect 22540 65548 22596 65550
rect 22988 69580 23044 69636
rect 22764 65996 22820 66052
rect 22428 64764 22484 64820
rect 23772 74508 23828 74564
rect 24220 74060 24276 74116
rect 23436 72492 23492 72548
rect 23212 70140 23268 70196
rect 23548 70700 23604 70756
rect 23100 69132 23156 69188
rect 23772 72658 23828 72660
rect 23772 72606 23774 72658
rect 23774 72606 23826 72658
rect 23826 72606 23828 72658
rect 23772 72604 23828 72606
rect 23772 71090 23828 71092
rect 23772 71038 23774 71090
rect 23774 71038 23826 71090
rect 23826 71038 23828 71090
rect 23772 71036 23828 71038
rect 27916 78652 27972 78708
rect 25116 77980 25172 78036
rect 24668 75068 24724 75124
rect 24892 75740 24948 75796
rect 27804 77756 27860 77812
rect 27692 77532 27748 77588
rect 27468 77420 27524 77476
rect 24668 74898 24724 74900
rect 24668 74846 24670 74898
rect 24670 74846 24722 74898
rect 24722 74846 24724 74898
rect 24668 74844 24724 74846
rect 24444 73388 24500 73444
rect 24780 73724 24836 73780
rect 24332 72716 24388 72772
rect 23996 72380 24052 72436
rect 24444 72546 24500 72548
rect 24444 72494 24446 72546
rect 24446 72494 24498 72546
rect 24498 72494 24500 72546
rect 24444 72492 24500 72494
rect 24892 71932 24948 71988
rect 23660 70588 23716 70644
rect 23436 67842 23492 67844
rect 23436 67790 23438 67842
rect 23438 67790 23490 67842
rect 23490 67790 23492 67842
rect 23436 67788 23492 67790
rect 23884 70588 23940 70644
rect 24332 70700 24388 70756
rect 24332 70194 24388 70196
rect 24332 70142 24334 70194
rect 24334 70142 24386 70194
rect 24386 70142 24388 70194
rect 24332 70140 24388 70142
rect 24108 68348 24164 68404
rect 23212 67564 23268 67620
rect 23548 66444 23604 66500
rect 23100 64818 23156 64820
rect 23100 64766 23102 64818
rect 23102 64766 23154 64818
rect 23154 64766 23156 64818
rect 23100 64764 23156 64766
rect 22428 64482 22484 64484
rect 22428 64430 22430 64482
rect 22430 64430 22482 64482
rect 22482 64430 22484 64482
rect 22428 64428 22484 64430
rect 22988 64204 23044 64260
rect 22204 63922 22260 63924
rect 22204 63870 22206 63922
rect 22206 63870 22258 63922
rect 22258 63870 22260 63922
rect 22204 63868 22260 63870
rect 22988 63868 23044 63924
rect 22316 63532 22372 63588
rect 21756 62860 21812 62916
rect 21084 62748 21140 62804
rect 21532 62578 21588 62580
rect 21532 62526 21534 62578
rect 21534 62526 21586 62578
rect 21586 62526 21588 62578
rect 21532 62524 21588 62526
rect 22876 63362 22932 63364
rect 22876 63310 22878 63362
rect 22878 63310 22930 63362
rect 22930 63310 22932 63362
rect 22876 63308 22932 63310
rect 22764 63084 22820 63140
rect 22092 62748 22148 62804
rect 22092 62524 22148 62580
rect 22204 62466 22260 62468
rect 22204 62414 22206 62466
rect 22206 62414 22258 62466
rect 22258 62414 22260 62466
rect 22204 62412 22260 62414
rect 21980 62188 22036 62244
rect 21756 61682 21812 61684
rect 21756 61630 21758 61682
rect 21758 61630 21810 61682
rect 21810 61630 21812 61682
rect 21756 61628 21812 61630
rect 21308 61292 21364 61348
rect 22204 61740 22260 61796
rect 20524 60172 20580 60228
rect 20860 60396 20916 60452
rect 20860 59724 20916 59780
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 22540 62748 22596 62804
rect 22316 61010 22372 61012
rect 22316 60958 22318 61010
rect 22318 60958 22370 61010
rect 22370 60958 22372 61010
rect 22316 60956 22372 60958
rect 22652 62188 22708 62244
rect 23436 65996 23492 66052
rect 23324 64764 23380 64820
rect 23884 67842 23940 67844
rect 23884 67790 23886 67842
rect 23886 67790 23938 67842
rect 23938 67790 23940 67842
rect 23884 67788 23940 67790
rect 24108 67452 24164 67508
rect 23772 65324 23828 65380
rect 23996 66946 24052 66948
rect 23996 66894 23998 66946
rect 23998 66894 24050 66946
rect 24050 66894 24052 66946
rect 23996 66892 24052 66894
rect 23884 64988 23940 65044
rect 23436 64204 23492 64260
rect 23548 64876 23604 64932
rect 23436 63980 23492 64036
rect 23212 63420 23268 63476
rect 23324 63532 23380 63588
rect 22652 61346 22708 61348
rect 22652 61294 22654 61346
rect 22654 61294 22706 61346
rect 22706 61294 22708 61346
rect 22652 61292 22708 61294
rect 23100 61180 23156 61236
rect 22204 60396 22260 60452
rect 23772 64876 23828 64932
rect 23996 64818 24052 64820
rect 23996 64766 23998 64818
rect 23998 64766 24050 64818
rect 24050 64766 24052 64818
rect 23996 64764 24052 64766
rect 23884 64706 23940 64708
rect 23884 64654 23886 64706
rect 23886 64654 23938 64706
rect 23938 64654 23940 64706
rect 23884 64652 23940 64654
rect 24220 67228 24276 67284
rect 24332 69580 24388 69636
rect 24444 68460 24500 68516
rect 24444 67900 24500 67956
rect 24556 67618 24612 67620
rect 24556 67566 24558 67618
rect 24558 67566 24610 67618
rect 24610 67566 24612 67618
rect 24556 67564 24612 67566
rect 24444 67452 24500 67508
rect 24220 65490 24276 65492
rect 24220 65438 24222 65490
rect 24222 65438 24274 65490
rect 24274 65438 24276 65490
rect 24220 65436 24276 65438
rect 24444 65266 24500 65268
rect 24444 65214 24446 65266
rect 24446 65214 24498 65266
rect 24498 65214 24500 65266
rect 24444 65212 24500 65214
rect 24332 64428 24388 64484
rect 24108 64146 24164 64148
rect 24108 64094 24110 64146
rect 24110 64094 24162 64146
rect 24162 64094 24164 64146
rect 24108 64092 24164 64094
rect 23884 63868 23940 63924
rect 23660 63644 23716 63700
rect 23660 63250 23716 63252
rect 23660 63198 23662 63250
rect 23662 63198 23714 63250
rect 23714 63198 23716 63250
rect 23660 63196 23716 63198
rect 23660 62636 23716 62692
rect 23548 61964 23604 62020
rect 23436 61180 23492 61236
rect 24220 63698 24276 63700
rect 24220 63646 24222 63698
rect 24222 63646 24274 63698
rect 24274 63646 24276 63698
rect 24220 63644 24276 63646
rect 23884 63308 23940 63364
rect 24108 63420 24164 63476
rect 23772 61964 23828 62020
rect 23772 61628 23828 61684
rect 23212 60674 23268 60676
rect 23212 60622 23214 60674
rect 23214 60622 23266 60674
rect 23266 60622 23268 60674
rect 23212 60620 23268 60622
rect 23212 60114 23268 60116
rect 23212 60062 23214 60114
rect 23214 60062 23266 60114
rect 23266 60062 23268 60114
rect 23212 60060 23268 60062
rect 24332 63362 24388 63364
rect 24332 63310 24334 63362
rect 24334 63310 24386 63362
rect 24386 63310 24388 63362
rect 24332 63308 24388 63310
rect 24220 63196 24276 63252
rect 24220 62636 24276 62692
rect 24556 63420 24612 63476
rect 24892 70252 24948 70308
rect 24892 69916 24948 69972
rect 24780 68348 24836 68404
rect 24780 67900 24836 67956
rect 25116 73052 25172 73108
rect 27132 76076 27188 76132
rect 25788 75458 25844 75460
rect 25788 75406 25790 75458
rect 25790 75406 25842 75458
rect 25842 75406 25844 75458
rect 25788 75404 25844 75406
rect 27020 74956 27076 75012
rect 25676 74786 25732 74788
rect 25676 74734 25678 74786
rect 25678 74734 25730 74786
rect 25730 74734 25732 74786
rect 25676 74732 25732 74734
rect 25340 71372 25396 71428
rect 25564 74620 25620 74676
rect 25228 71202 25284 71204
rect 25228 71150 25230 71202
rect 25230 71150 25282 71202
rect 25282 71150 25284 71202
rect 25228 71148 25284 71150
rect 26348 73612 26404 73668
rect 26684 73612 26740 73668
rect 26124 73500 26180 73556
rect 25676 73218 25732 73220
rect 25676 73166 25678 73218
rect 25678 73166 25730 73218
rect 25730 73166 25732 73218
rect 25676 73164 25732 73166
rect 25788 72322 25844 72324
rect 25788 72270 25790 72322
rect 25790 72270 25842 72322
rect 25842 72270 25844 72322
rect 25788 72268 25844 72270
rect 25676 71762 25732 71764
rect 25676 71710 25678 71762
rect 25678 71710 25730 71762
rect 25730 71710 25732 71762
rect 25676 71708 25732 71710
rect 25452 70866 25508 70868
rect 25452 70814 25454 70866
rect 25454 70814 25506 70866
rect 25506 70814 25508 70866
rect 25452 70812 25508 70814
rect 25116 70476 25172 70532
rect 25116 70140 25172 70196
rect 25116 69244 25172 69300
rect 25340 69132 25396 69188
rect 26572 72156 26628 72212
rect 26348 71820 26404 71876
rect 26236 71484 26292 71540
rect 26572 71484 26628 71540
rect 25452 68124 25508 68180
rect 26012 70700 26068 70756
rect 25676 70082 25732 70084
rect 25676 70030 25678 70082
rect 25678 70030 25730 70082
rect 25730 70030 25732 70082
rect 25676 70028 25732 70030
rect 26460 69916 26516 69972
rect 26012 69692 26068 69748
rect 25676 68796 25732 68852
rect 26460 69468 26516 69524
rect 26572 70028 26628 70084
rect 26124 69410 26180 69412
rect 26124 69358 26126 69410
rect 26126 69358 26178 69410
rect 26178 69358 26180 69410
rect 26124 69356 26180 69358
rect 26012 69020 26068 69076
rect 26124 68908 26180 68964
rect 26348 68796 26404 68852
rect 25900 68348 25956 68404
rect 26012 68572 26068 68628
rect 25564 68012 25620 68068
rect 26236 68626 26292 68628
rect 26236 68574 26238 68626
rect 26238 68574 26290 68626
rect 26290 68574 26292 68626
rect 26236 68572 26292 68574
rect 25788 67452 25844 67508
rect 25340 66556 25396 66612
rect 25452 66892 25508 66948
rect 24892 65884 24948 65940
rect 25452 66220 25508 66276
rect 24892 65548 24948 65604
rect 25116 65660 25172 65716
rect 24780 63532 24836 63588
rect 24892 65324 24948 65380
rect 25116 65100 25172 65156
rect 24892 64204 24948 64260
rect 24220 61682 24276 61684
rect 24220 61630 24222 61682
rect 24222 61630 24274 61682
rect 24274 61630 24276 61682
rect 24220 61628 24276 61630
rect 24668 62636 24724 62692
rect 25116 64706 25172 64708
rect 25116 64654 25118 64706
rect 25118 64654 25170 64706
rect 25170 64654 25172 64706
rect 25116 64652 25172 64654
rect 25564 66162 25620 66164
rect 25564 66110 25566 66162
rect 25566 66110 25618 66162
rect 25618 66110 25620 66162
rect 25564 66108 25620 66110
rect 25676 64764 25732 64820
rect 25452 64540 25508 64596
rect 25676 64594 25732 64596
rect 25676 64542 25678 64594
rect 25678 64542 25730 64594
rect 25730 64542 25732 64594
rect 25676 64540 25732 64542
rect 26348 67340 26404 67396
rect 26236 67228 26292 67284
rect 26124 67170 26180 67172
rect 26124 67118 26126 67170
rect 26126 67118 26178 67170
rect 26178 67118 26180 67170
rect 26124 67116 26180 67118
rect 26236 66556 26292 66612
rect 26908 71538 26964 71540
rect 26908 71486 26910 71538
rect 26910 71486 26962 71538
rect 26962 71486 26964 71538
rect 26908 71484 26964 71486
rect 27020 71372 27076 71428
rect 27132 74060 27188 74116
rect 27356 73500 27412 73556
rect 27244 73276 27300 73332
rect 27244 70812 27300 70868
rect 26796 70028 26852 70084
rect 26572 68908 26628 68964
rect 26796 68908 26852 68964
rect 27916 77644 27972 77700
rect 27804 73218 27860 73220
rect 27804 73166 27806 73218
rect 27806 73166 27858 73218
rect 27858 73166 27860 73218
rect 27804 73164 27860 73166
rect 28028 77532 28084 77588
rect 28588 77532 28644 77588
rect 28140 76466 28196 76468
rect 28140 76414 28142 76466
rect 28142 76414 28194 76466
rect 28194 76414 28196 76466
rect 28140 76412 28196 76414
rect 28700 76412 28756 76468
rect 28364 75852 28420 75908
rect 28364 75068 28420 75124
rect 31836 76860 31892 76916
rect 31724 76636 31780 76692
rect 29820 75794 29876 75796
rect 29820 75742 29822 75794
rect 29822 75742 29874 75794
rect 29874 75742 29876 75794
rect 29820 75740 29876 75742
rect 29036 75292 29092 75348
rect 28588 72492 28644 72548
rect 28924 73836 28980 73892
rect 28812 73500 28868 73556
rect 28812 73164 28868 73220
rect 28812 72546 28868 72548
rect 28812 72494 28814 72546
rect 28814 72494 28866 72546
rect 28866 72494 28868 72546
rect 28812 72492 28868 72494
rect 28252 72156 28308 72212
rect 27580 71762 27636 71764
rect 27580 71710 27582 71762
rect 27582 71710 27634 71762
rect 27634 71710 27636 71762
rect 27580 71708 27636 71710
rect 27468 71260 27524 71316
rect 27580 70476 27636 70532
rect 27580 69804 27636 69860
rect 27692 70588 27748 70644
rect 27132 69410 27188 69412
rect 27132 69358 27134 69410
rect 27134 69358 27186 69410
rect 27186 69358 27188 69410
rect 27132 69356 27188 69358
rect 26796 67452 26852 67508
rect 26796 67058 26852 67060
rect 26796 67006 26798 67058
rect 26798 67006 26850 67058
rect 26850 67006 26852 67058
rect 26796 67004 26852 67006
rect 26012 65996 26068 66052
rect 27356 67900 27412 67956
rect 27468 67788 27524 67844
rect 27132 67170 27188 67172
rect 27132 67118 27134 67170
rect 27134 67118 27186 67170
rect 27186 67118 27188 67170
rect 27132 67116 27188 67118
rect 27020 66332 27076 66388
rect 27356 66780 27412 66836
rect 26908 66274 26964 66276
rect 26908 66222 26910 66274
rect 26910 66222 26962 66274
rect 26962 66222 26964 66274
rect 26908 66220 26964 66222
rect 27132 66274 27188 66276
rect 27132 66222 27134 66274
rect 27134 66222 27186 66274
rect 27186 66222 27188 66274
rect 27132 66220 27188 66222
rect 26012 65490 26068 65492
rect 26012 65438 26014 65490
rect 26014 65438 26066 65490
rect 26066 65438 26068 65490
rect 26012 65436 26068 65438
rect 26460 65490 26516 65492
rect 26460 65438 26462 65490
rect 26462 65438 26514 65490
rect 26514 65438 26516 65490
rect 26460 65436 26516 65438
rect 25900 64876 25956 64932
rect 26348 65324 26404 65380
rect 26684 65324 26740 65380
rect 26348 65100 26404 65156
rect 26684 64706 26740 64708
rect 26684 64654 26686 64706
rect 26686 64654 26738 64706
rect 26738 64654 26740 64706
rect 26684 64652 26740 64654
rect 25788 64034 25844 64036
rect 25788 63982 25790 64034
rect 25790 63982 25842 64034
rect 25842 63982 25844 64034
rect 25788 63980 25844 63982
rect 25116 63644 25172 63700
rect 25116 63084 25172 63140
rect 26572 64092 26628 64148
rect 27356 65660 27412 65716
rect 27468 65548 27524 65604
rect 27020 65436 27076 65492
rect 27580 65436 27636 65492
rect 28028 69410 28084 69412
rect 28028 69358 28030 69410
rect 28030 69358 28082 69410
rect 28082 69358 28084 69410
rect 28028 69356 28084 69358
rect 27804 68236 27860 68292
rect 28028 68796 28084 68852
rect 29148 73442 29204 73444
rect 29148 73390 29150 73442
rect 29150 73390 29202 73442
rect 29202 73390 29204 73442
rect 29148 73388 29204 73390
rect 29036 72716 29092 72772
rect 30492 75740 30548 75796
rect 30380 74844 30436 74900
rect 29932 74172 29988 74228
rect 29372 73330 29428 73332
rect 29372 73278 29374 73330
rect 29374 73278 29426 73330
rect 29426 73278 29428 73330
rect 29372 73276 29428 73278
rect 28812 71932 28868 71988
rect 28364 69580 28420 69636
rect 28588 69580 28644 69636
rect 28588 69410 28644 69412
rect 28588 69358 28590 69410
rect 28590 69358 28642 69410
rect 28642 69358 28644 69410
rect 28588 69356 28644 69358
rect 28364 69020 28420 69076
rect 28476 69244 28532 69300
rect 28252 68796 28308 68852
rect 28028 67452 28084 67508
rect 27916 66892 27972 66948
rect 27804 65996 27860 66052
rect 28252 67116 28308 67172
rect 28364 66332 28420 66388
rect 28028 65660 28084 65716
rect 26908 64988 26964 65044
rect 27020 64930 27076 64932
rect 27020 64878 27022 64930
rect 27022 64878 27074 64930
rect 27074 64878 27076 64930
rect 27020 64876 27076 64878
rect 27468 64988 27524 65044
rect 27132 64092 27188 64148
rect 26460 63868 26516 63924
rect 25900 63756 25956 63812
rect 25900 62636 25956 62692
rect 26348 62636 26404 62692
rect 26908 63922 26964 63924
rect 26908 63870 26910 63922
rect 26910 63870 26962 63922
rect 26962 63870 26964 63922
rect 26908 63868 26964 63870
rect 27132 63868 27188 63924
rect 26684 63756 26740 63812
rect 28140 65436 28196 65492
rect 28364 64876 28420 64932
rect 28252 64818 28308 64820
rect 28252 64766 28254 64818
rect 28254 64766 28306 64818
rect 28306 64766 28308 64818
rect 28252 64764 28308 64766
rect 28252 63980 28308 64036
rect 28812 68908 28868 68964
rect 28700 68514 28756 68516
rect 28700 68462 28702 68514
rect 28702 68462 28754 68514
rect 28754 68462 28756 68514
rect 28700 68460 28756 68462
rect 28812 67954 28868 67956
rect 28812 67902 28814 67954
rect 28814 67902 28866 67954
rect 28866 67902 28868 67954
rect 28812 67900 28868 67902
rect 28588 67170 28644 67172
rect 28588 67118 28590 67170
rect 28590 67118 28642 67170
rect 28642 67118 28644 67170
rect 28588 67116 28644 67118
rect 28812 67004 28868 67060
rect 28700 66892 28756 66948
rect 28588 65660 28644 65716
rect 27580 63084 27636 63140
rect 26796 62914 26852 62916
rect 26796 62862 26798 62914
rect 26798 62862 26850 62914
rect 26850 62862 26852 62914
rect 26796 62860 26852 62862
rect 27692 62860 27748 62916
rect 28252 63084 28308 63140
rect 29820 73164 29876 73220
rect 29708 72828 29764 72884
rect 29820 72604 29876 72660
rect 29148 71762 29204 71764
rect 29148 71710 29150 71762
rect 29150 71710 29202 71762
rect 29202 71710 29204 71762
rect 29148 71708 29204 71710
rect 29372 70924 29428 70980
rect 29484 71596 29540 71652
rect 29372 70476 29428 70532
rect 29036 69356 29092 69412
rect 29148 68572 29204 68628
rect 29148 68124 29204 68180
rect 29596 71484 29652 71540
rect 29708 71372 29764 71428
rect 29596 71202 29652 71204
rect 29596 71150 29598 71202
rect 29598 71150 29650 71202
rect 29650 71150 29652 71202
rect 29596 71148 29652 71150
rect 29708 71036 29764 71092
rect 30044 74508 30100 74564
rect 30268 74508 30324 74564
rect 30268 74114 30324 74116
rect 30268 74062 30270 74114
rect 30270 74062 30322 74114
rect 30322 74062 30324 74114
rect 30268 74060 30324 74062
rect 30268 72828 30324 72884
rect 31836 76578 31892 76580
rect 31836 76526 31838 76578
rect 31838 76526 31890 76578
rect 31890 76526 31892 76578
rect 31836 76524 31892 76526
rect 30940 76300 30996 76356
rect 30604 75292 30660 75348
rect 30828 74898 30884 74900
rect 30828 74846 30830 74898
rect 30830 74846 30882 74898
rect 30882 74846 30884 74898
rect 30828 74844 30884 74846
rect 30604 74284 30660 74340
rect 30492 73500 30548 73556
rect 30492 73052 30548 73108
rect 30940 73276 30996 73332
rect 30604 72940 30660 72996
rect 30492 72658 30548 72660
rect 30492 72606 30494 72658
rect 30494 72606 30546 72658
rect 30546 72606 30548 72658
rect 30492 72604 30548 72606
rect 30268 72156 30324 72212
rect 29596 70306 29652 70308
rect 29596 70254 29598 70306
rect 29598 70254 29650 70306
rect 29650 70254 29652 70306
rect 29596 70252 29652 70254
rect 29820 70306 29876 70308
rect 29820 70254 29822 70306
rect 29822 70254 29874 70306
rect 29874 70254 29876 70306
rect 29820 70252 29876 70254
rect 30044 71484 30100 71540
rect 30156 71260 30212 71316
rect 30380 70978 30436 70980
rect 30380 70926 30382 70978
rect 30382 70926 30434 70978
rect 30434 70926 30436 70978
rect 30380 70924 30436 70926
rect 30380 70700 30436 70756
rect 30940 72716 30996 72772
rect 30604 72268 30660 72324
rect 30828 72380 30884 72436
rect 30604 71762 30660 71764
rect 30604 71710 30606 71762
rect 30606 71710 30658 71762
rect 30658 71710 30660 71762
rect 30604 71708 30660 71710
rect 30492 70252 30548 70308
rect 30044 70028 30100 70084
rect 30044 69804 30100 69860
rect 30156 69468 30212 69524
rect 29708 68796 29764 68852
rect 30268 69356 30324 69412
rect 30044 69298 30100 69300
rect 30044 69246 30046 69298
rect 30046 69246 30098 69298
rect 30098 69246 30100 69298
rect 30044 69244 30100 69246
rect 29932 69186 29988 69188
rect 29932 69134 29934 69186
rect 29934 69134 29986 69186
rect 29986 69134 29988 69186
rect 29932 69132 29988 69134
rect 30044 69020 30100 69076
rect 29932 68908 29988 68964
rect 29596 68066 29652 68068
rect 29596 68014 29598 68066
rect 29598 68014 29650 68066
rect 29650 68014 29652 68066
rect 29596 68012 29652 68014
rect 29372 67900 29428 67956
rect 29820 67900 29876 67956
rect 29148 67116 29204 67172
rect 29372 67170 29428 67172
rect 29372 67118 29374 67170
rect 29374 67118 29426 67170
rect 29426 67118 29428 67170
rect 29372 67116 29428 67118
rect 28924 66668 28980 66724
rect 29596 67058 29652 67060
rect 29596 67006 29598 67058
rect 29598 67006 29650 67058
rect 29650 67006 29652 67058
rect 29596 67004 29652 67006
rect 29708 66892 29764 66948
rect 29596 66220 29652 66276
rect 29372 65772 29428 65828
rect 29932 67730 29988 67732
rect 29932 67678 29934 67730
rect 29934 67678 29986 67730
rect 29986 67678 29988 67730
rect 29932 67676 29988 67678
rect 29708 65660 29764 65716
rect 28812 65100 28868 65156
rect 28924 65324 28980 65380
rect 29932 65772 29988 65828
rect 29484 65324 29540 65380
rect 29820 64818 29876 64820
rect 29820 64766 29822 64818
rect 29822 64766 29874 64818
rect 29874 64766 29876 64818
rect 29820 64764 29876 64766
rect 28924 64146 28980 64148
rect 28924 64094 28926 64146
rect 28926 64094 28978 64146
rect 28978 64094 28980 64146
rect 28924 64092 28980 64094
rect 28812 63084 28868 63140
rect 29932 63138 29988 63140
rect 29932 63086 29934 63138
rect 29934 63086 29986 63138
rect 29986 63086 29988 63138
rect 29932 63084 29988 63086
rect 28364 62524 28420 62580
rect 28476 63026 28532 63028
rect 28476 62974 28478 63026
rect 28478 62974 28530 63026
rect 28530 62974 28532 63026
rect 28476 62972 28532 62974
rect 25340 62188 25396 62244
rect 24892 61964 24948 62020
rect 25116 61964 25172 62020
rect 24556 61628 24612 61684
rect 25004 61852 25060 61908
rect 21308 59388 21364 59444
rect 19516 58940 19572 58996
rect 19628 58828 19684 58884
rect 19180 57932 19236 57988
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 18620 56588 18676 56644
rect 19516 57148 19572 57204
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 21868 55356 21924 55412
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 25900 61682 25956 61684
rect 25900 61630 25902 61682
rect 25902 61630 25954 61682
rect 25954 61630 25956 61682
rect 25900 61628 25956 61630
rect 28028 61404 28084 61460
rect 29596 63026 29652 63028
rect 29596 62974 29598 63026
rect 29598 62974 29650 63026
rect 29650 62974 29652 63026
rect 29596 62972 29652 62974
rect 28812 62578 28868 62580
rect 28812 62526 28814 62578
rect 28814 62526 28866 62578
rect 28866 62526 28868 62578
rect 28812 62524 28868 62526
rect 29708 61740 29764 61796
rect 29820 61404 29876 61460
rect 30828 69298 30884 69300
rect 30828 69246 30830 69298
rect 30830 69246 30882 69298
rect 30882 69246 30884 69298
rect 30828 69244 30884 69246
rect 30716 68908 30772 68964
rect 30716 68572 30772 68628
rect 30604 67900 30660 67956
rect 32060 76748 32116 76804
rect 36764 76748 36820 76804
rect 33404 76524 33460 76580
rect 34636 76578 34692 76580
rect 34636 76526 34638 76578
rect 34638 76526 34690 76578
rect 34690 76526 34692 76578
rect 34636 76524 34692 76526
rect 35980 76578 36036 76580
rect 35980 76526 35982 76578
rect 35982 76526 36034 76578
rect 36034 76526 36036 76578
rect 35980 76524 36036 76526
rect 35532 76412 35588 76468
rect 32396 76188 32452 76244
rect 31276 75740 31332 75796
rect 31388 75628 31444 75684
rect 31948 75682 32004 75684
rect 31948 75630 31950 75682
rect 31950 75630 32002 75682
rect 32002 75630 32004 75682
rect 31948 75628 32004 75630
rect 31164 74396 31220 74452
rect 31612 74732 31668 74788
rect 31388 74226 31444 74228
rect 31388 74174 31390 74226
rect 31390 74174 31442 74226
rect 31442 74174 31444 74226
rect 31388 74172 31444 74174
rect 31500 73330 31556 73332
rect 31500 73278 31502 73330
rect 31502 73278 31554 73330
rect 31554 73278 31556 73330
rect 31500 73276 31556 73278
rect 31164 72940 31220 72996
rect 31164 72604 31220 72660
rect 31052 70924 31108 70980
rect 31052 70252 31108 70308
rect 31948 74508 32004 74564
rect 32956 75570 33012 75572
rect 32956 75518 32958 75570
rect 32958 75518 33010 75570
rect 33010 75518 33012 75570
rect 32956 75516 33012 75518
rect 32172 74732 32228 74788
rect 32284 74172 32340 74228
rect 31836 72716 31892 72772
rect 32060 72658 32116 72660
rect 32060 72606 32062 72658
rect 32062 72606 32114 72658
rect 32114 72606 32116 72658
rect 32060 72604 32116 72606
rect 31836 72268 31892 72324
rect 31724 71932 31780 71988
rect 31276 70028 31332 70084
rect 31164 69804 31220 69860
rect 31052 69468 31108 69524
rect 31388 68684 31444 68740
rect 31724 70700 31780 70756
rect 32732 74284 32788 74340
rect 33068 74956 33124 75012
rect 32508 74114 32564 74116
rect 32508 74062 32510 74114
rect 32510 74062 32562 74114
rect 32562 74062 32564 74114
rect 32508 74060 32564 74062
rect 32732 73164 32788 73220
rect 31836 69580 31892 69636
rect 32284 73052 32340 73108
rect 32620 72716 32676 72772
rect 32396 71986 32452 71988
rect 32396 71934 32398 71986
rect 32398 71934 32450 71986
rect 32450 71934 32452 71986
rect 32396 71932 32452 71934
rect 33180 74844 33236 74900
rect 33404 74396 33460 74452
rect 34636 76300 34692 76356
rect 33740 75964 33796 76020
rect 33740 75740 33796 75796
rect 34188 75682 34244 75684
rect 34188 75630 34190 75682
rect 34190 75630 34242 75682
rect 34242 75630 34244 75682
rect 34188 75628 34244 75630
rect 34524 74898 34580 74900
rect 34524 74846 34526 74898
rect 34526 74846 34578 74898
rect 34578 74846 34580 74898
rect 34524 74844 34580 74846
rect 33852 74674 33908 74676
rect 33852 74622 33854 74674
rect 33854 74622 33906 74674
rect 33906 74622 33908 74674
rect 33852 74620 33908 74622
rect 33628 74396 33684 74452
rect 34076 74060 34132 74116
rect 34412 74114 34468 74116
rect 34412 74062 34414 74114
rect 34414 74062 34466 74114
rect 34466 74062 34468 74114
rect 34412 74060 34468 74062
rect 33180 73890 33236 73892
rect 33180 73838 33182 73890
rect 33182 73838 33234 73890
rect 33234 73838 33236 73890
rect 33180 73836 33236 73838
rect 32844 73052 32900 73108
rect 31724 69356 31780 69412
rect 31836 69020 31892 69076
rect 31724 68908 31780 68964
rect 31500 68572 31556 68628
rect 31612 68684 31668 68740
rect 31388 68514 31444 68516
rect 31388 68462 31390 68514
rect 31390 68462 31442 68514
rect 31442 68462 31444 68514
rect 31388 68460 31444 68462
rect 31836 68684 31892 68740
rect 31388 67900 31444 67956
rect 32396 70476 32452 70532
rect 32284 70194 32340 70196
rect 32284 70142 32286 70194
rect 32286 70142 32338 70194
rect 32338 70142 32340 70194
rect 32284 70140 32340 70142
rect 32060 70028 32116 70084
rect 32172 69916 32228 69972
rect 32396 70028 32452 70084
rect 32284 68626 32340 68628
rect 32284 68574 32286 68626
rect 32286 68574 32338 68626
rect 32338 68574 32340 68626
rect 32284 68572 32340 68574
rect 32620 69804 32676 69860
rect 32956 71484 33012 71540
rect 33516 73276 33572 73332
rect 33740 73052 33796 73108
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 33964 73164 34020 73220
rect 35756 76188 35812 76244
rect 36540 76300 36596 76356
rect 38668 77756 38724 77812
rect 37772 76524 37828 76580
rect 37884 77644 37940 77700
rect 36764 76300 36820 76356
rect 35644 75628 35700 75684
rect 36092 75570 36148 75572
rect 36092 75518 36094 75570
rect 36094 75518 36146 75570
rect 36146 75518 36148 75570
rect 36092 75516 36148 75518
rect 35420 74844 35476 74900
rect 34860 74732 34916 74788
rect 34860 74508 34916 74564
rect 34748 72940 34804 72996
rect 33852 72322 33908 72324
rect 33852 72270 33854 72322
rect 33854 72270 33906 72322
rect 33906 72270 33908 72322
rect 33852 72268 33908 72270
rect 34748 72268 34804 72324
rect 33852 71874 33908 71876
rect 33852 71822 33854 71874
rect 33854 71822 33906 71874
rect 33906 71822 33908 71874
rect 33852 71820 33908 71822
rect 33404 71148 33460 71204
rect 33404 70978 33460 70980
rect 33404 70926 33406 70978
rect 33406 70926 33458 70978
rect 33458 70926 33460 70978
rect 33404 70924 33460 70926
rect 32844 70364 32900 70420
rect 33292 70700 33348 70756
rect 32732 69634 32788 69636
rect 32732 69582 32734 69634
rect 32734 69582 32786 69634
rect 32786 69582 32788 69634
rect 32732 69580 32788 69582
rect 32620 69244 32676 69300
rect 32508 69132 32564 69188
rect 32508 68796 32564 68852
rect 32620 68460 32676 68516
rect 31948 67564 32004 67620
rect 31388 67116 31444 67172
rect 31276 67058 31332 67060
rect 31276 67006 31278 67058
rect 31278 67006 31330 67058
rect 31330 67006 31332 67058
rect 31276 67004 31332 67006
rect 31276 66668 31332 66724
rect 31948 66668 32004 66724
rect 30604 65772 30660 65828
rect 30492 65714 30548 65716
rect 30492 65662 30494 65714
rect 30494 65662 30546 65714
rect 30546 65662 30548 65714
rect 30492 65660 30548 65662
rect 30380 65548 30436 65604
rect 30268 65490 30324 65492
rect 30268 65438 30270 65490
rect 30270 65438 30322 65490
rect 30322 65438 30324 65490
rect 30268 65436 30324 65438
rect 31052 65714 31108 65716
rect 31052 65662 31054 65714
rect 31054 65662 31106 65714
rect 31106 65662 31108 65714
rect 31052 65660 31108 65662
rect 31276 65548 31332 65604
rect 31500 65324 31556 65380
rect 30044 61180 30100 61236
rect 30380 62860 30436 62916
rect 30380 60284 30436 60340
rect 28476 57036 28532 57092
rect 28812 56588 28868 56644
rect 25116 55132 25172 55188
rect 27804 56252 27860 56308
rect 25116 54908 25172 54964
rect 26012 54908 26068 54964
rect 21868 49980 21924 50036
rect 23212 49980 23268 50036
rect 19516 48524 19572 48580
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 17612 36706 17668 36708
rect 17612 36654 17614 36706
rect 17614 36654 17666 36706
rect 17666 36654 17668 36706
rect 17612 36652 17668 36654
rect 17612 36204 17668 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 17500 6748 17556 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18620 5964 18676 6020
rect 19628 6018 19684 6020
rect 19628 5966 19630 6018
rect 19630 5966 19682 6018
rect 19682 5966 19684 6018
rect 19628 5964 19684 5966
rect 18172 5794 18228 5796
rect 18172 5742 18174 5794
rect 18174 5742 18226 5794
rect 18226 5742 18228 5794
rect 18172 5740 18228 5742
rect 18844 5740 18900 5796
rect 16716 5292 16772 5348
rect 18844 5068 18900 5124
rect 15372 4508 15428 4564
rect 11676 3612 11732 3668
rect 12236 3666 12292 3668
rect 12236 3614 12238 3666
rect 12238 3614 12290 3666
rect 12290 3614 12292 3666
rect 12236 3612 12292 3614
rect 16604 4450 16660 4452
rect 16604 4398 16606 4450
rect 16606 4398 16658 4450
rect 16658 4398 16660 4450
rect 16604 4396 16660 4398
rect 17500 4396 17556 4452
rect 26012 5180 26068 5236
rect 22204 5122 22260 5124
rect 22204 5070 22206 5122
rect 22206 5070 22258 5122
rect 22258 5070 22260 5122
rect 22204 5068 22260 5070
rect 23436 5122 23492 5124
rect 23436 5070 23438 5122
rect 23438 5070 23490 5122
rect 23490 5070 23492 5122
rect 23436 5068 23492 5070
rect 26796 5068 26852 5124
rect 24668 4898 24724 4900
rect 24668 4846 24670 4898
rect 24670 4846 24722 4898
rect 24722 4846 24724 4898
rect 24668 4844 24724 4846
rect 26012 4844 26068 4900
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 15148 3612 15204 3668
rect 16044 3666 16100 3668
rect 16044 3614 16046 3666
rect 16046 3614 16098 3666
rect 16098 3614 16100 3666
rect 16044 3612 16100 3614
rect 16380 3612 16436 3668
rect 19964 4450 20020 4452
rect 19964 4398 19966 4450
rect 19966 4398 20018 4450
rect 20018 4398 20020 4450
rect 19964 4396 20020 4398
rect 21420 4396 21476 4452
rect 18172 3666 18228 3668
rect 18172 3614 18174 3666
rect 18174 3614 18226 3666
rect 18226 3614 18228 3666
rect 18172 3612 18228 3614
rect 21084 3612 21140 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 25788 3612 25844 3668
rect 28812 55468 28868 55524
rect 29596 55468 29652 55524
rect 32508 67618 32564 67620
rect 32508 67566 32510 67618
rect 32510 67566 32562 67618
rect 32562 67566 32564 67618
rect 32508 67564 32564 67566
rect 32844 68908 32900 68964
rect 32956 68850 33012 68852
rect 32956 68798 32958 68850
rect 32958 68798 33010 68850
rect 33010 68798 33012 68850
rect 32956 68796 33012 68798
rect 32844 68738 32900 68740
rect 32844 68686 32846 68738
rect 32846 68686 32898 68738
rect 32898 68686 32900 68738
rect 32844 68684 32900 68686
rect 32396 67170 32452 67172
rect 32396 67118 32398 67170
rect 32398 67118 32450 67170
rect 32450 67118 32452 67170
rect 32396 67116 32452 67118
rect 32844 67170 32900 67172
rect 32844 67118 32846 67170
rect 32846 67118 32898 67170
rect 32898 67118 32900 67170
rect 32844 67116 32900 67118
rect 33740 70418 33796 70420
rect 33740 70366 33742 70418
rect 33742 70366 33794 70418
rect 33794 70366 33796 70418
rect 33740 70364 33796 70366
rect 33516 69916 33572 69972
rect 33516 69634 33572 69636
rect 33516 69582 33518 69634
rect 33518 69582 33570 69634
rect 33570 69582 33572 69634
rect 33516 69580 33572 69582
rect 33404 69410 33460 69412
rect 33404 69358 33406 69410
rect 33406 69358 33458 69410
rect 33458 69358 33460 69410
rect 33404 69356 33460 69358
rect 33516 69244 33572 69300
rect 34076 69580 34132 69636
rect 34076 69410 34132 69412
rect 34076 69358 34078 69410
rect 34078 69358 34130 69410
rect 34130 69358 34132 69410
rect 34076 69356 34132 69358
rect 33852 68796 33908 68852
rect 33964 69132 34020 69188
rect 33516 68738 33572 68740
rect 33516 68686 33518 68738
rect 33518 68686 33570 68738
rect 33570 68686 33572 68738
rect 33516 68684 33572 68686
rect 34188 68124 34244 68180
rect 33964 67730 34020 67732
rect 33964 67678 33966 67730
rect 33966 67678 34018 67730
rect 34018 67678 34020 67730
rect 33964 67676 34020 67678
rect 33516 66892 33572 66948
rect 34636 70978 34692 70980
rect 34636 70926 34638 70978
rect 34638 70926 34690 70978
rect 34690 70926 34692 70978
rect 34636 70924 34692 70926
rect 34636 70082 34692 70084
rect 34636 70030 34638 70082
rect 34638 70030 34690 70082
rect 34690 70030 34692 70082
rect 34636 70028 34692 70030
rect 37548 76076 37604 76132
rect 36988 75068 37044 75124
rect 36764 74786 36820 74788
rect 36764 74734 36766 74786
rect 36766 74734 36818 74786
rect 36818 74734 36820 74786
rect 36764 74732 36820 74734
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 36092 74396 36148 74452
rect 34972 74060 35028 74116
rect 35196 74172 35252 74228
rect 35980 74114 36036 74116
rect 35980 74062 35982 74114
rect 35982 74062 36034 74114
rect 36034 74062 36036 74114
rect 35980 74060 36036 74062
rect 35644 73724 35700 73780
rect 35084 73052 35140 73108
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35644 72716 35700 72772
rect 35980 72828 36036 72884
rect 35980 72434 36036 72436
rect 35980 72382 35982 72434
rect 35982 72382 36034 72434
rect 36034 72382 36036 72434
rect 35980 72380 36036 72382
rect 35084 72322 35140 72324
rect 35084 72270 35086 72322
rect 35086 72270 35138 72322
rect 35138 72270 35140 72322
rect 35084 72268 35140 72270
rect 35084 71874 35140 71876
rect 35084 71822 35086 71874
rect 35086 71822 35138 71874
rect 35138 71822 35140 71874
rect 35084 71820 35140 71822
rect 35532 71874 35588 71876
rect 35532 71822 35534 71874
rect 35534 71822 35586 71874
rect 35586 71822 35588 71874
rect 35532 71820 35588 71822
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 71148 35252 71204
rect 35980 71148 36036 71204
rect 35532 71090 35588 71092
rect 35532 71038 35534 71090
rect 35534 71038 35586 71090
rect 35586 71038 35588 71090
rect 35532 71036 35588 71038
rect 34860 70364 34916 70420
rect 35084 70306 35140 70308
rect 35084 70254 35086 70306
rect 35086 70254 35138 70306
rect 35138 70254 35140 70306
rect 35084 70252 35140 70254
rect 35532 70028 35588 70084
rect 35756 70140 35812 70196
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35308 69580 35364 69636
rect 35532 68796 35588 68852
rect 34524 68684 34580 68740
rect 34412 68514 34468 68516
rect 34412 68462 34414 68514
rect 34414 68462 34466 68514
rect 34466 68462 34468 68514
rect 34412 68460 34468 68462
rect 34412 67788 34468 67844
rect 35308 68348 35364 68404
rect 34860 68124 34916 68180
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 34412 67618 34468 67620
rect 34412 67566 34414 67618
rect 34414 67566 34466 67618
rect 34466 67566 34468 67618
rect 34412 67564 34468 67566
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 36316 74620 36372 74676
rect 36540 74284 36596 74340
rect 36428 73724 36484 73780
rect 36316 73052 36372 73108
rect 36428 72658 36484 72660
rect 36428 72606 36430 72658
rect 36430 72606 36482 72658
rect 36482 72606 36484 72658
rect 36428 72604 36484 72606
rect 36428 72156 36484 72212
rect 35980 67452 36036 67508
rect 36316 72044 36372 72100
rect 35532 66444 35588 66500
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 34300 63196 34356 63252
rect 33292 61964 33348 62020
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 33180 56812 33236 56868
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 29932 55074 29988 55076
rect 29932 55022 29934 55074
rect 29934 55022 29986 55074
rect 29986 55022 29988 55074
rect 29932 55020 29988 55022
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 36876 73442 36932 73444
rect 36876 73390 36878 73442
rect 36878 73390 36930 73442
rect 36930 73390 36932 73442
rect 36876 73388 36932 73390
rect 36876 71986 36932 71988
rect 36876 71934 36878 71986
rect 36878 71934 36930 71986
rect 36930 71934 36932 71986
rect 36876 71932 36932 71934
rect 36876 71596 36932 71652
rect 36428 70418 36484 70420
rect 36428 70366 36430 70418
rect 36430 70366 36482 70418
rect 36482 70366 36484 70418
rect 36428 70364 36484 70366
rect 37212 74786 37268 74788
rect 37212 74734 37214 74786
rect 37214 74734 37266 74786
rect 37266 74734 37268 74786
rect 37212 74732 37268 74734
rect 37436 74172 37492 74228
rect 38332 76860 38388 76916
rect 38220 75852 38276 75908
rect 37660 74786 37716 74788
rect 37660 74734 37662 74786
rect 37662 74734 37714 74786
rect 37714 74734 37716 74786
rect 37660 74732 37716 74734
rect 37100 70924 37156 70980
rect 37884 74226 37940 74228
rect 37884 74174 37886 74226
rect 37886 74174 37938 74226
rect 37938 74174 37940 74226
rect 37884 74172 37940 74174
rect 37324 73554 37380 73556
rect 37324 73502 37326 73554
rect 37326 73502 37378 73554
rect 37378 73502 37380 73554
rect 37324 73500 37380 73502
rect 38556 75122 38612 75124
rect 38556 75070 38558 75122
rect 38558 75070 38610 75122
rect 38610 75070 38612 75122
rect 38556 75068 38612 75070
rect 40124 77532 40180 77588
rect 39900 76690 39956 76692
rect 39900 76638 39902 76690
rect 39902 76638 39954 76690
rect 39954 76638 39956 76690
rect 39900 76636 39956 76638
rect 39004 76578 39060 76580
rect 39004 76526 39006 76578
rect 39006 76526 39058 76578
rect 39058 76526 39060 76578
rect 39004 76524 39060 76526
rect 38780 76300 38836 76356
rect 40908 77420 40964 77476
rect 42140 76524 42196 76580
rect 43372 76578 43428 76580
rect 43372 76526 43374 76578
rect 43374 76526 43426 76578
rect 43426 76526 43428 76578
rect 43372 76524 43428 76526
rect 48860 77980 48916 78036
rect 46508 76524 46564 76580
rect 47628 76578 47684 76580
rect 47628 76526 47630 76578
rect 47630 76526 47682 76578
rect 47682 76526 47684 76578
rect 47628 76524 47684 76526
rect 48748 76578 48804 76580
rect 48748 76526 48750 76578
rect 48750 76526 48802 76578
rect 48802 76526 48804 76578
rect 48748 76524 48804 76526
rect 39452 75628 39508 75684
rect 39228 75292 39284 75348
rect 38668 73836 38724 73892
rect 37772 72044 37828 72100
rect 37772 71762 37828 71764
rect 37772 71710 37774 71762
rect 37774 71710 37826 71762
rect 37826 71710 37828 71762
rect 37772 71708 37828 71710
rect 37772 70588 37828 70644
rect 37212 70476 37268 70532
rect 36988 70194 37044 70196
rect 36988 70142 36990 70194
rect 36990 70142 37042 70194
rect 37042 70142 37044 70194
rect 36988 70140 37044 70142
rect 37324 70194 37380 70196
rect 37324 70142 37326 70194
rect 37326 70142 37378 70194
rect 37378 70142 37380 70194
rect 37324 70140 37380 70142
rect 37884 68684 37940 68740
rect 36204 68460 36260 68516
rect 38780 73164 38836 73220
rect 38332 72546 38388 72548
rect 38332 72494 38334 72546
rect 38334 72494 38386 72546
rect 38386 72494 38388 72546
rect 38332 72492 38388 72494
rect 38780 72546 38836 72548
rect 38780 72494 38782 72546
rect 38782 72494 38834 72546
rect 38834 72494 38836 72546
rect 38780 72492 38836 72494
rect 38668 72156 38724 72212
rect 38332 63756 38388 63812
rect 38108 60172 38164 60228
rect 39228 73164 39284 73220
rect 39564 73218 39620 73220
rect 39564 73166 39566 73218
rect 39566 73166 39618 73218
rect 39618 73166 39620 73218
rect 39564 73164 39620 73166
rect 41468 74786 41524 74788
rect 41468 74734 41470 74786
rect 41470 74734 41522 74786
rect 41522 74734 41524 74786
rect 41468 74732 41524 74734
rect 41356 72044 41412 72100
rect 42364 73724 42420 73780
rect 46620 72380 46676 72436
rect 41916 71708 41972 71764
rect 40796 68796 40852 68852
rect 39116 66780 39172 66836
rect 38668 58156 38724 58212
rect 40348 66332 40404 66388
rect 38668 57596 38724 57652
rect 40012 57596 40068 57652
rect 36092 51996 36148 52052
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 32620 41916 32676 41972
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34300 5234 34356 5236
rect 34300 5182 34302 5234
rect 34302 5182 34354 5234
rect 34354 5182 34356 5234
rect 34300 5180 34356 5182
rect 28028 5068 28084 5124
rect 32060 5122 32116 5124
rect 32060 5070 32062 5122
rect 32062 5070 32114 5122
rect 32114 5070 32116 5122
rect 32060 5068 32116 5070
rect 33292 5122 33348 5124
rect 33292 5070 33294 5122
rect 33294 5070 33346 5122
rect 33346 5070 33348 5122
rect 33292 5068 33348 5070
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34748 5234 34804 5236
rect 34748 5182 34750 5234
rect 34750 5182 34802 5234
rect 34802 5182 34804 5234
rect 34748 5180 34804 5182
rect 40348 54684 40404 54740
rect 47852 59276 47908 59332
rect 40348 53788 40404 53844
rect 41244 53788 41300 53844
rect 34412 5068 34468 5124
rect 34972 5122 35028 5124
rect 34972 5070 34974 5122
rect 34974 5070 35026 5122
rect 35026 5070 35028 5122
rect 34972 5068 35028 5070
rect 39452 5122 39508 5124
rect 39452 5070 39454 5122
rect 39454 5070 39506 5122
rect 39506 5070 39508 5122
rect 39452 5068 39508 5070
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 29596 4450 29652 4452
rect 29596 4398 29598 4450
rect 29598 4398 29650 4450
rect 29650 4398 29652 4450
rect 29596 4396 29652 4398
rect 30716 4396 30772 4452
rect 28364 4338 28420 4340
rect 28364 4286 28366 4338
rect 28366 4286 28418 4338
rect 28418 4286 28420 4338
rect 28364 4284 28420 4286
rect 29260 4338 29316 4340
rect 29260 4286 29262 4338
rect 29262 4286 29314 4338
rect 29314 4286 29316 4338
rect 29260 4284 29316 4286
rect 26684 3666 26740 3668
rect 26684 3614 26686 3666
rect 26686 3614 26738 3666
rect 26738 3614 26740 3666
rect 26684 3612 26740 3614
rect 30492 3612 30548 3668
rect 31388 3666 31444 3668
rect 31388 3614 31390 3666
rect 31390 3614 31442 3666
rect 31442 3614 31444 3666
rect 31388 3612 31444 3614
rect 35308 4396 35364 4452
rect 38332 4450 38388 4452
rect 38332 4398 38334 4450
rect 38334 4398 38386 4450
rect 38386 4398 38388 4450
rect 38332 4396 38388 4398
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35196 3612 35252 3668
rect 35756 3666 35812 3668
rect 35756 3614 35758 3666
rect 35758 3614 35810 3666
rect 35810 3614 35812 3666
rect 35756 3612 35812 3614
rect 41020 4396 41076 4452
rect 38668 3500 38724 3556
rect 39900 3612 39956 3668
rect 41020 3554 41076 3556
rect 41020 3502 41022 3554
rect 41022 3502 41074 3554
rect 41074 3502 41076 3554
rect 41020 3500 41076 3502
rect 46844 5292 46900 5348
rect 47740 5292 47796 5348
rect 47180 5122 47236 5124
rect 47180 5070 47182 5122
rect 47182 5070 47234 5122
rect 47234 5070 47236 5122
rect 47180 5068 47236 5070
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50876 76524 50932 76580
rect 51548 76578 51604 76580
rect 51548 76526 51550 76578
rect 51550 76526 51602 76578
rect 51602 76526 51604 76578
rect 51548 76524 51604 76526
rect 52668 76578 52724 76580
rect 52668 76526 52670 76578
rect 52670 76526 52722 76578
rect 52722 76526 52724 76578
rect 52668 76524 52724 76526
rect 59948 76524 60004 76580
rect 61628 76578 61684 76580
rect 61628 76526 61630 76578
rect 61630 76526 61682 76578
rect 61682 76526 61684 76578
rect 61628 76524 61684 76526
rect 67788 76748 67844 76804
rect 68348 76748 68404 76804
rect 69580 76748 69636 76804
rect 63980 76524 64036 76580
rect 65548 76578 65604 76580
rect 65548 76526 65550 76578
rect 65550 76526 65602 76578
rect 65602 76526 65604 76578
rect 65548 76524 65604 76526
rect 74956 77308 75012 77364
rect 72716 76524 72772 76580
rect 72940 76636 72996 76692
rect 55244 75516 55300 75572
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 56476 75570 56532 75572
rect 56476 75518 56478 75570
rect 56478 75518 56530 75570
rect 56530 75518 56532 75570
rect 56476 75516 56532 75518
rect 60620 74620 60676 74676
rect 73948 76578 74004 76580
rect 73948 76526 73950 76578
rect 73950 76526 74002 76578
rect 74002 76526 74004 76578
rect 73948 76524 74004 76526
rect 68572 76188 68628 76244
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 64540 74060 64596 74116
rect 55356 72828 55412 72884
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50428 71820 50484 71876
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 77308 55020 77364 55076
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 48860 50316 48916 50372
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 48860 49756 48916 49812
rect 49532 49756 49588 49812
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 49532 6076 49588 6132
rect 51212 6130 51268 6132
rect 51212 6078 51214 6130
rect 51214 6078 51266 6130
rect 51266 6078 51268 6130
rect 51212 6076 51268 6078
rect 52220 6076 52276 6132
rect 52892 5852 52948 5908
rect 47964 5122 48020 5124
rect 47964 5070 47966 5122
rect 47966 5070 48018 5122
rect 48018 5070 48020 5122
rect 47964 5068 48020 5070
rect 51212 5068 51268 5124
rect 47852 4508 47908 4564
rect 43484 4450 43540 4452
rect 43484 4398 43486 4450
rect 43486 4398 43538 4450
rect 43538 4398 43540 4450
rect 43484 4396 43540 4398
rect 41692 3666 41748 3668
rect 41692 3614 41694 3666
rect 41694 3614 41746 3666
rect 41746 3614 41748 3666
rect 41692 3612 41748 3614
rect 41244 3500 41300 3556
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50764 4562 50820 4564
rect 50764 4510 50766 4562
rect 50766 4510 50818 4562
rect 50818 4510 50820 4562
rect 50764 4508 50820 4510
rect 51772 5068 51828 5124
rect 51996 5068 52052 5124
rect 51772 4508 51828 4564
rect 48300 4396 48356 4452
rect 49532 4450 49588 4452
rect 49532 4398 49534 4450
rect 49534 4398 49586 4450
rect 49586 4398 49588 4450
rect 49532 4396 49588 4398
rect 49868 4450 49924 4452
rect 49868 4398 49870 4450
rect 49870 4398 49922 4450
rect 49922 4398 49924 4450
rect 49868 4396 49924 4398
rect 50540 4396 50596 4452
rect 52332 5122 52388 5124
rect 52332 5070 52334 5122
rect 52334 5070 52386 5122
rect 52386 5070 52388 5122
rect 52332 5068 52388 5070
rect 52780 4396 52836 4452
rect 53340 5852 53396 5908
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 53004 5068 53060 5124
rect 52332 4226 52388 4228
rect 52332 4174 52334 4226
rect 52334 4174 52386 4226
rect 52386 4174 52388 4226
rect 52332 4172 52388 4174
rect 53452 4338 53508 4340
rect 53452 4286 53454 4338
rect 53454 4286 53506 4338
rect 53506 4286 53508 4338
rect 53452 4284 53508 4286
rect 54012 4338 54068 4340
rect 54012 4286 54014 4338
rect 54014 4286 54066 4338
rect 54066 4286 54068 4338
rect 54012 4284 54068 4286
rect 54012 3612 54068 3668
rect 51660 3554 51716 3556
rect 51660 3502 51662 3554
rect 51662 3502 51714 3554
rect 51714 3502 51716 3554
rect 51660 3500 51716 3502
rect 52780 3554 52836 3556
rect 52780 3502 52782 3554
rect 52782 3502 52834 3554
rect 52834 3502 52836 3554
rect 52780 3500 52836 3502
rect 53340 3554 53396 3556
rect 53340 3502 53342 3554
rect 53342 3502 53394 3554
rect 53394 3502 53396 3554
rect 53340 3500 53396 3502
rect 45612 3388 45668 3444
rect 44604 3276 44660 3332
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 54908 4450 54964 4452
rect 54908 4398 54910 4450
rect 54910 4398 54962 4450
rect 54962 4398 54964 4450
rect 54908 4396 54964 4398
rect 55244 4450 55300 4452
rect 55244 4398 55246 4450
rect 55246 4398 55298 4450
rect 55298 4398 55300 4450
rect 55244 4396 55300 4398
rect 58268 4450 58324 4452
rect 58268 4398 58270 4450
rect 58270 4398 58322 4450
rect 58322 4398 58324 4450
rect 58268 4396 58324 4398
rect 64540 4396 64596 4452
rect 57932 4172 57988 4228
rect 58604 4284 58660 4340
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 58716 3612 58772 3668
rect 59276 3666 59332 3668
rect 59276 3614 59278 3666
rect 59278 3614 59330 3666
rect 59330 3614 59332 3666
rect 59276 3612 59332 3614
rect 63420 3612 63476 3668
rect 66220 4450 66276 4452
rect 66220 4398 66222 4450
rect 66222 4398 66274 4450
rect 66274 4398 66276 4450
rect 66220 4396 66276 4398
rect 68460 4396 68516 4452
rect 65324 4284 65380 4340
rect 65884 4338 65940 4340
rect 65884 4286 65886 4338
rect 65886 4286 65938 4338
rect 65938 4286 65940 4338
rect 65884 4284 65940 4286
rect 65212 3666 65268 3668
rect 65212 3614 65214 3666
rect 65214 3614 65266 3666
rect 65266 3614 65268 3666
rect 65212 3612 65268 3614
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65324 3500 65380 3556
rect 68124 3612 68180 3668
rect 74396 4338 74452 4340
rect 74396 4286 74398 4338
rect 74398 4286 74450 4338
rect 74450 4286 74452 4338
rect 74396 4284 74452 4286
rect 75180 4338 75236 4340
rect 75180 4286 75182 4338
rect 75182 4286 75234 4338
rect 75234 4286 75236 4338
rect 75180 4284 75236 4286
rect 76076 4226 76132 4228
rect 76076 4174 76078 4226
rect 76078 4174 76130 4226
rect 76130 4174 76132 4226
rect 76076 4172 76132 4174
rect 69132 3666 69188 3668
rect 69132 3614 69134 3666
rect 69134 3614 69186 3666
rect 69186 3614 69188 3666
rect 69132 3612 69188 3614
rect 72828 3612 72884 3668
rect 72604 3554 72660 3556
rect 72604 3502 72606 3554
rect 72606 3502 72658 3554
rect 72658 3502 72660 3554
rect 72604 3500 72660 3502
rect 73724 3666 73780 3668
rect 73724 3614 73726 3666
rect 73726 3614 73778 3666
rect 73778 3614 73780 3666
rect 73724 3612 73780 3614
rect 73276 3554 73332 3556
rect 73276 3502 73278 3554
rect 73278 3502 73330 3554
rect 73330 3502 73332 3554
rect 73276 3500 73332 3502
rect 77420 36204 77476 36260
rect 77420 4284 77476 4340
rect 77308 3500 77364 3556
rect 77532 4172 77588 4228
<< metal3 >>
rect 3042 79884 3052 79940
rect 3108 79884 14364 79940
rect 14420 79884 14430 79940
rect 2380 79660 14476 79716
rect 14532 79660 28812 79716
rect 28868 79660 28878 79716
rect 2380 79044 2436 79660
rect 10882 79548 10892 79604
rect 10948 79548 28364 79604
rect 28420 79548 28430 79604
rect 4946 79436 4956 79492
rect 5012 79436 17948 79492
rect 18004 79436 18014 79492
rect 8306 79324 8316 79380
rect 8372 79324 15148 79380
rect 15204 79324 15214 79380
rect 8866 79212 8876 79268
rect 8932 79212 21532 79268
rect 21588 79212 21598 79268
rect 4498 79100 4508 79156
rect 4564 79100 18396 79156
rect 18452 79100 18462 79156
rect 2370 78988 2380 79044
rect 2436 78988 2446 79044
rect 4162 78988 4172 79044
rect 4228 78988 18732 79044
rect 18788 78988 18798 79044
rect 5842 78876 5852 78932
rect 5908 78876 17388 78932
rect 17444 78876 17454 78932
rect 2034 78764 2044 78820
rect 2100 78764 15932 78820
rect 15988 78764 15998 78820
rect 3826 78652 3836 78708
rect 3892 78652 27916 78708
rect 27972 78652 27982 78708
rect 2930 78540 2940 78596
rect 2996 78540 20412 78596
rect 20468 78540 20478 78596
rect 4834 78428 4844 78484
rect 4900 78428 24556 78484
rect 24612 78428 24622 78484
rect 3378 78316 3388 78372
rect 3444 78316 22988 78372
rect 23044 78316 23054 78372
rect 7634 78204 7644 78260
rect 7700 78204 17612 78260
rect 17668 78204 17678 78260
rect 6738 78092 6748 78148
rect 6804 78092 20188 78148
rect 20244 78092 20254 78148
rect 4946 77980 4956 78036
rect 5012 77980 19068 78036
rect 19124 77980 19134 78036
rect 25106 77980 25116 78036
rect 25172 77980 48860 78036
rect 48916 77980 48926 78036
rect 2706 77868 2716 77924
rect 2772 77868 14588 77924
rect 14644 77868 14654 77924
rect 2482 77756 2492 77812
rect 2548 77756 3388 77812
rect 4274 77756 4284 77812
rect 4340 77756 8428 77812
rect 8484 77756 8494 77812
rect 9090 77756 9100 77812
rect 9156 77756 27804 77812
rect 27860 77756 38668 77812
rect 38724 77756 38734 77812
rect 3332 77700 3388 77756
rect 3332 77644 7084 77700
rect 7140 77644 7150 77700
rect 7298 77644 7308 77700
rect 7364 77644 20188 77700
rect 27906 77644 27916 77700
rect 27972 77644 37884 77700
rect 37940 77644 37950 77700
rect 20132 77588 20188 77644
rect 4610 77532 4620 77588
rect 4676 77532 7644 77588
rect 7700 77532 12124 77588
rect 12180 77532 12190 77588
rect 20132 77532 27692 77588
rect 27748 77532 27758 77588
rect 28018 77532 28028 77588
rect 28084 77532 28588 77588
rect 28644 77532 40124 77588
rect 40180 77532 40190 77588
rect 4050 77420 4060 77476
rect 4116 77420 10220 77476
rect 10276 77420 10286 77476
rect 12226 77420 12236 77476
rect 12292 77420 27468 77476
rect 27524 77420 40908 77476
rect 40964 77420 40974 77476
rect 2146 77308 2156 77364
rect 2212 77308 4732 77364
rect 4788 77308 4956 77364
rect 5012 77308 5022 77364
rect 5180 77308 11452 77364
rect 11508 77308 13804 77364
rect 13860 77308 13870 77364
rect 14028 77308 23548 77364
rect 23604 77308 23614 77364
rect 24210 77308 24220 77364
rect 24276 77308 74956 77364
rect 75012 77308 75022 77364
rect 5180 77252 5236 77308
rect 14028 77252 14084 77308
rect 3490 77196 3500 77252
rect 3556 77196 5236 77252
rect 9650 77196 9660 77252
rect 9716 77196 14084 77252
rect 3266 76860 3276 76916
rect 3332 76860 9996 76916
rect 10052 76860 12012 76916
rect 12068 76860 12078 76916
rect 31826 76860 31836 76916
rect 31892 76860 38332 76916
rect 38388 76860 38398 76916
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 3266 76748 3276 76804
rect 3332 76748 6636 76804
rect 6692 76748 6702 76804
rect 32050 76748 32060 76804
rect 32116 76748 33292 76804
rect 33348 76748 36764 76804
rect 36820 76748 36830 76804
rect 67778 76748 67788 76804
rect 67844 76748 68348 76804
rect 68404 76748 69580 76804
rect 69636 76748 69646 76804
rect 3938 76636 3948 76692
rect 4004 76636 11564 76692
rect 11620 76636 11630 76692
rect 12114 76636 12124 76692
rect 12180 76636 31724 76692
rect 31780 76636 39900 76692
rect 39956 76636 39966 76692
rect 43652 76636 72940 76692
rect 72996 76636 73006 76692
rect 3490 76524 3500 76580
rect 3556 76524 6524 76580
rect 6580 76524 6590 76580
rect 8418 76524 8428 76580
rect 8484 76524 18844 76580
rect 18900 76524 18910 76580
rect 20626 76524 20636 76580
rect 20692 76524 31836 76580
rect 31892 76524 31902 76580
rect 33394 76524 33404 76580
rect 33460 76524 34636 76580
rect 34692 76524 35980 76580
rect 36036 76524 36046 76580
rect 37762 76524 37772 76580
rect 37828 76524 39004 76580
rect 39060 76524 39070 76580
rect 42130 76524 42140 76580
rect 42196 76524 43372 76580
rect 43428 76524 43438 76580
rect 43652 76468 43708 76636
rect 46498 76524 46508 76580
rect 46564 76524 47628 76580
rect 47684 76524 48748 76580
rect 48804 76524 48814 76580
rect 50866 76524 50876 76580
rect 50932 76524 51548 76580
rect 51604 76524 52668 76580
rect 52724 76524 52734 76580
rect 59938 76524 59948 76580
rect 60004 76524 61628 76580
rect 61684 76524 61694 76580
rect 63970 76524 63980 76580
rect 64036 76524 65548 76580
rect 65604 76524 65614 76580
rect 72706 76524 72716 76580
rect 72772 76524 73948 76580
rect 74004 76524 74014 76580
rect 2034 76412 2044 76468
rect 2100 76412 4396 76468
rect 4452 76412 4462 76468
rect 6290 76412 6300 76468
rect 6356 76412 7308 76468
rect 7364 76412 7374 76468
rect 16706 76412 16716 76468
rect 16772 76412 20300 76468
rect 20356 76412 20366 76468
rect 22306 76412 22316 76468
rect 22372 76412 24332 76468
rect 24388 76412 28140 76468
rect 28196 76412 28700 76468
rect 28756 76412 28766 76468
rect 35522 76412 35532 76468
rect 35588 76412 43708 76468
rect 3490 76300 3500 76356
rect 3556 76300 4508 76356
rect 4564 76300 4574 76356
rect 6626 76300 6636 76356
rect 6692 76300 13580 76356
rect 13636 76300 13646 76356
rect 15092 76300 18508 76356
rect 18564 76300 18574 76356
rect 21382 76300 21420 76356
rect 21476 76300 21486 76356
rect 30930 76300 30940 76356
rect 30996 76300 34636 76356
rect 34692 76300 36540 76356
rect 36596 76300 36606 76356
rect 36754 76300 36764 76356
rect 36820 76300 38780 76356
rect 38836 76300 38846 76356
rect 15092 76244 15148 76300
rect 3602 76188 3612 76244
rect 3668 76188 4340 76244
rect 4610 76188 4620 76244
rect 4676 76188 5628 76244
rect 5684 76188 5694 76244
rect 6290 76188 6300 76244
rect 6356 76188 10668 76244
rect 10724 76188 10734 76244
rect 10994 76188 11004 76244
rect 11060 76188 15148 76244
rect 15922 76188 15932 76244
rect 15988 76188 30604 76244
rect 30660 76188 30670 76244
rect 32386 76188 32396 76244
rect 32452 76188 35588 76244
rect 35746 76188 35756 76244
rect 35812 76188 68572 76244
rect 68628 76188 68638 76244
rect 3378 75964 3388 76020
rect 3444 75964 3612 76020
rect 3668 75964 3836 76020
rect 3892 75964 3902 76020
rect 4284 75908 4340 76188
rect 35532 76132 35588 76188
rect 6738 76076 6748 76132
rect 6804 76076 9996 76132
rect 10052 76076 10062 76132
rect 11554 76076 11564 76132
rect 11620 76076 18060 76132
rect 18116 76076 18126 76132
rect 20132 76076 27132 76132
rect 27188 76076 27198 76132
rect 35532 76076 37548 76132
rect 37604 76076 37614 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 20132 76020 20188 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 9874 75964 9884 76020
rect 9940 75964 10892 76020
rect 10948 75964 10958 76020
rect 13794 75964 13804 76020
rect 13860 75964 15484 76020
rect 15540 75964 20188 76020
rect 26852 75964 33740 76020
rect 33796 75964 33806 76020
rect 2006 75852 2044 75908
rect 2100 75852 2110 75908
rect 4284 75852 5404 75908
rect 5460 75852 5470 75908
rect 5954 75852 5964 75908
rect 6020 75852 6972 75908
rect 7028 75852 10668 75908
rect 10724 75852 10734 75908
rect 12114 75852 12124 75908
rect 12180 75852 12348 75908
rect 12404 75852 12414 75908
rect 13458 75852 13468 75908
rect 13524 75852 13916 75908
rect 13972 75852 18620 75908
rect 18676 75852 18686 75908
rect 26852 75796 26908 75964
rect 28354 75852 28364 75908
rect 28420 75852 38220 75908
rect 38276 75852 38286 75908
rect 3714 75740 3724 75796
rect 3780 75740 7980 75796
rect 8036 75740 8046 75796
rect 8194 75740 8204 75796
rect 8260 75740 9212 75796
rect 9268 75740 9278 75796
rect 10546 75740 10556 75796
rect 10612 75740 12908 75796
rect 12964 75740 14140 75796
rect 14196 75740 14206 75796
rect 16818 75740 16828 75796
rect 16884 75740 23156 75796
rect 24882 75740 24892 75796
rect 24948 75740 26908 75796
rect 29810 75740 29820 75796
rect 29876 75740 30492 75796
rect 30548 75740 31276 75796
rect 31332 75740 31342 75796
rect 33730 75740 33740 75796
rect 33796 75740 38668 75796
rect 23100 75684 23156 75740
rect 38612 75684 38668 75740
rect 4162 75628 4172 75684
rect 4228 75628 4508 75684
rect 4564 75628 4574 75684
rect 6850 75628 6860 75684
rect 6916 75628 8988 75684
rect 9044 75628 10108 75684
rect 10164 75628 14028 75684
rect 14084 75628 16940 75684
rect 16996 75628 17500 75684
rect 17556 75628 17566 75684
rect 20290 75628 20300 75684
rect 20356 75628 22316 75684
rect 22372 75628 22382 75684
rect 23100 75628 26124 75684
rect 26180 75628 26190 75684
rect 31378 75628 31388 75684
rect 31444 75628 31948 75684
rect 32004 75628 32014 75684
rect 34178 75628 34188 75684
rect 34244 75628 35644 75684
rect 35700 75628 35710 75684
rect 38612 75628 39452 75684
rect 39508 75628 39518 75684
rect 2594 75516 2604 75572
rect 2660 75516 3724 75572
rect 3780 75516 3948 75572
rect 4004 75516 4014 75572
rect 4386 75516 4396 75572
rect 4452 75516 4462 75572
rect 4722 75516 4732 75572
rect 4788 75516 7196 75572
rect 7252 75516 7262 75572
rect 7522 75516 7532 75572
rect 7588 75516 13692 75572
rect 13748 75516 13758 75572
rect 17714 75516 17724 75572
rect 17780 75516 19404 75572
rect 19460 75516 19470 75572
rect 32946 75516 32956 75572
rect 33012 75516 36092 75572
rect 36148 75516 36158 75572
rect 55234 75516 55244 75572
rect 55300 75516 56476 75572
rect 56532 75516 56542 75572
rect 4396 75460 4452 75516
rect 2034 75404 2044 75460
rect 2100 75404 2828 75460
rect 2884 75404 2894 75460
rect 3826 75404 3836 75460
rect 3892 75404 3902 75460
rect 4050 75404 4060 75460
rect 4116 75404 4452 75460
rect 4834 75404 4844 75460
rect 4900 75404 7532 75460
rect 7588 75404 7598 75460
rect 8754 75404 8764 75460
rect 8820 75404 11340 75460
rect 11396 75404 13468 75460
rect 13524 75404 13534 75460
rect 13794 75404 13804 75460
rect 13860 75404 18396 75460
rect 18452 75404 18462 75460
rect 22978 75404 22988 75460
rect 23044 75404 25788 75460
rect 25844 75404 25854 75460
rect 3042 75180 3052 75236
rect 3108 75180 3500 75236
rect 3556 75180 3566 75236
rect 3836 75012 3892 75404
rect 8194 75292 8204 75348
rect 8260 75292 10780 75348
rect 10836 75292 13412 75348
rect 13682 75292 13692 75348
rect 13748 75292 18172 75348
rect 18228 75292 18238 75348
rect 29026 75292 29036 75348
rect 29092 75292 30604 75348
rect 30660 75292 39228 75348
rect 39284 75292 39294 75348
rect 13356 75124 13412 75292
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 5730 75068 5740 75124
rect 5796 75068 13132 75124
rect 13188 75068 13198 75124
rect 13356 75068 17724 75124
rect 17780 75068 17790 75124
rect 24658 75068 24668 75124
rect 24724 75068 28364 75124
rect 28420 75068 28430 75124
rect 29586 75068 29596 75124
rect 29652 75068 33628 75124
rect 33684 75068 33694 75124
rect 36978 75068 36988 75124
rect 37044 75068 38556 75124
rect 38612 75068 38622 75124
rect 3836 74956 4060 75012
rect 4116 74956 4126 75012
rect 5170 74956 5180 75012
rect 5236 74956 7756 75012
rect 7812 74956 8652 75012
rect 8708 74956 9884 75012
rect 9940 74956 9950 75012
rect 13010 74956 13020 75012
rect 13076 74956 15148 75012
rect 15204 74956 15214 75012
rect 16034 74956 16044 75012
rect 16100 74956 18732 75012
rect 18788 74956 18798 75012
rect 20132 74956 27020 75012
rect 27076 74956 27086 75012
rect 30594 74956 30604 75012
rect 30660 74956 33068 75012
rect 33124 74956 38668 75012
rect 20132 74900 20188 74956
rect 3332 74844 4956 74900
rect 5012 74844 5022 74900
rect 5282 74844 5292 74900
rect 5348 74844 8764 74900
rect 8820 74844 8830 74900
rect 8978 74844 8988 74900
rect 9044 74844 9772 74900
rect 9828 74844 11116 74900
rect 11172 74844 11182 74900
rect 12674 74844 12684 74900
rect 12740 74844 20188 74900
rect 24658 74844 24668 74900
rect 24724 74844 30380 74900
rect 30436 74844 30446 74900
rect 30818 74844 30828 74900
rect 30884 74844 33180 74900
rect 33236 74844 34524 74900
rect 34580 74844 35420 74900
rect 35476 74844 35486 74900
rect 3332 74788 3388 74844
rect 38612 74788 38668 74956
rect 2594 74732 2604 74788
rect 2660 74732 3388 74788
rect 4162 74732 4172 74788
rect 4228 74732 4508 74788
rect 4564 74732 4574 74788
rect 10546 74732 10556 74788
rect 10612 74732 11788 74788
rect 11844 74732 11854 74788
rect 12012 74732 13356 74788
rect 13412 74732 13422 74788
rect 17490 74732 17500 74788
rect 17556 74732 22092 74788
rect 22148 74732 22158 74788
rect 25554 74732 25564 74788
rect 25620 74732 25676 74788
rect 25732 74732 25742 74788
rect 31602 74732 31612 74788
rect 31668 74732 32172 74788
rect 32228 74732 32238 74788
rect 34850 74732 34860 74788
rect 34916 74732 36764 74788
rect 36820 74732 37212 74788
rect 37268 74732 37660 74788
rect 37716 74732 37726 74788
rect 38612 74732 41468 74788
rect 41524 74732 41534 74788
rect 1586 74620 1596 74676
rect 1652 74620 2828 74676
rect 2884 74620 2894 74676
rect 3052 74620 6076 74676
rect 6132 74620 6142 74676
rect 7410 74620 7420 74676
rect 7476 74620 7532 74676
rect 7588 74620 7598 74676
rect 10294 74620 10332 74676
rect 10388 74620 10398 74676
rect 3052 74564 3108 74620
rect 12012 74564 12068 74732
rect 12450 74620 12460 74676
rect 12516 74620 13132 74676
rect 13188 74620 13198 74676
rect 13356 74620 21756 74676
rect 21812 74620 21822 74676
rect 25554 74620 25564 74676
rect 25620 74620 33852 74676
rect 33908 74620 36316 74676
rect 36372 74620 60620 74676
rect 60676 74620 60686 74676
rect 1250 74508 1260 74564
rect 1316 74508 3108 74564
rect 5506 74508 5516 74564
rect 5572 74508 12068 74564
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 13356 74452 13412 74620
rect 18386 74508 18396 74564
rect 18452 74508 18620 74564
rect 18676 74508 23772 74564
rect 23828 74508 30044 74564
rect 30100 74508 30110 74564
rect 30258 74508 30268 74564
rect 30324 74508 31948 74564
rect 32004 74508 32060 74564
rect 32116 74508 34860 74564
rect 34916 74508 34926 74564
rect 30044 74452 30100 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 36092 74452 36148 74620
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 7074 74396 7084 74452
rect 7140 74396 11788 74452
rect 11844 74396 13412 74452
rect 15138 74396 15148 74452
rect 15204 74396 20188 74452
rect 30044 74396 31164 74452
rect 31220 74396 33404 74452
rect 33460 74396 33628 74452
rect 33684 74396 33694 74452
rect 36082 74396 36092 74452
rect 36148 74396 36158 74452
rect 20132 74340 20188 74396
rect 33628 74340 33684 74396
rect 2370 74284 2380 74340
rect 2436 74284 3388 74340
rect 3444 74284 4060 74340
rect 4116 74284 4126 74340
rect 4946 74284 4956 74340
rect 5012 74284 8428 74340
rect 8484 74284 9660 74340
rect 9716 74284 9996 74340
rect 10052 74284 11452 74340
rect 11508 74284 11518 74340
rect 13458 74284 13468 74340
rect 13524 74284 16604 74340
rect 16660 74284 16670 74340
rect 20132 74284 30604 74340
rect 30660 74284 32732 74340
rect 32788 74284 32798 74340
rect 33628 74284 36540 74340
rect 36596 74284 36606 74340
rect 2818 74172 2828 74228
rect 2884 74172 5572 74228
rect 5730 74172 5740 74228
rect 5796 74172 8652 74228
rect 8708 74172 8718 74228
rect 11106 74172 11116 74228
rect 11172 74172 12684 74228
rect 12740 74172 12750 74228
rect 13346 74172 13356 74228
rect 13412 74172 20076 74228
rect 20132 74172 20142 74228
rect 29922 74172 29932 74228
rect 29988 74172 31388 74228
rect 31444 74172 31454 74228
rect 31602 74172 31612 74228
rect 31668 74172 32284 74228
rect 32340 74172 32564 74228
rect 35186 74172 35196 74228
rect 35252 74172 37436 74228
rect 37492 74172 37884 74228
rect 37940 74172 37950 74228
rect 5516 74116 5572 74172
rect 32508 74116 32564 74172
rect 2146 74060 2156 74116
rect 2212 74060 4396 74116
rect 4452 74060 4462 74116
rect 4722 74060 4732 74116
rect 4788 74060 5292 74116
rect 5348 74060 5358 74116
rect 5516 74060 7644 74116
rect 7700 74060 8204 74116
rect 8260 74060 8270 74116
rect 8372 74060 11004 74116
rect 11060 74060 11070 74116
rect 12002 74060 12012 74116
rect 12068 74060 14140 74116
rect 14196 74060 14206 74116
rect 15138 74060 15148 74116
rect 15204 74060 21532 74116
rect 21588 74060 21598 74116
rect 24210 74060 24220 74116
rect 24276 74060 26908 74116
rect 27122 74060 27132 74116
rect 27188 74060 30268 74116
rect 30324 74060 30334 74116
rect 32498 74060 32508 74116
rect 32564 74060 32574 74116
rect 34066 74060 34076 74116
rect 34132 74060 34412 74116
rect 34468 74060 34972 74116
rect 35028 74060 35980 74116
rect 36036 74060 64540 74116
rect 64596 74060 64606 74116
rect 8372 74004 8428 74060
rect 26852 74004 26908 74060
rect 3462 73948 3500 74004
rect 3556 73948 3566 74004
rect 3910 73948 3948 74004
rect 4004 73948 4014 74004
rect 6850 73948 6860 74004
rect 6916 73948 6972 74004
rect 7028 73948 7038 74004
rect 7186 73948 7196 74004
rect 7252 73948 7756 74004
rect 7812 73948 7822 74004
rect 7970 73948 7980 74004
rect 8036 73948 8092 74004
rect 8148 73948 8158 74004
rect 8316 73948 8428 74004
rect 9650 73948 9660 74004
rect 9716 73948 10108 74004
rect 10164 73948 10174 74004
rect 10434 73948 10444 74004
rect 10500 73948 11340 74004
rect 11396 73948 11406 74004
rect 11778 73948 11788 74004
rect 11844 73948 12124 74004
rect 12180 73948 12190 74004
rect 12786 73948 12796 74004
rect 12852 73948 16156 74004
rect 16212 73948 16222 74004
rect 21606 73948 21644 74004
rect 21700 73948 21710 74004
rect 22754 73948 22764 74004
rect 22820 73948 24836 74004
rect 26852 73948 29596 74004
rect 29652 73948 29662 74004
rect 31602 73948 31612 74004
rect 31668 73948 31678 74004
rect 33618 73948 33628 74004
rect 33684 73948 35252 74004
rect 8316 73892 8372 73948
rect 3826 73836 3836 73892
rect 3892 73836 5964 73892
rect 6020 73836 6030 73892
rect 6374 73836 6412 73892
rect 6468 73836 6478 73892
rect 6738 73836 6748 73892
rect 6804 73836 7196 73892
rect 7252 73836 7262 73892
rect 7420 73836 8372 73892
rect 8866 73836 8876 73892
rect 8932 73836 9436 73892
rect 9492 73836 9502 73892
rect 10434 73836 10444 73892
rect 10500 73836 11900 73892
rect 11956 73836 11966 73892
rect 14354 73836 14364 73892
rect 14420 73836 21868 73892
rect 21924 73836 21934 73892
rect 7420 73780 7476 73836
rect 24780 73780 24836 73948
rect 31612 73892 31668 73948
rect 35196 73892 35252 73948
rect 28914 73836 28924 73892
rect 28980 73836 31668 73892
rect 32946 73836 32956 73892
rect 33012 73836 33180 73892
rect 33236 73836 33246 73892
rect 35196 73836 38668 73892
rect 38724 73836 38734 73892
rect 4162 73724 4172 73780
rect 4228 73724 4844 73780
rect 4900 73724 4910 73780
rect 5282 73724 5292 73780
rect 5348 73724 7420 73780
rect 7476 73724 7486 73780
rect 8082 73724 8092 73780
rect 8148 73724 9996 73780
rect 10052 73724 10062 73780
rect 10210 73724 10220 73780
rect 10276 73724 10668 73780
rect 10724 73724 10734 73780
rect 24770 73724 24780 73780
rect 24836 73724 24846 73780
rect 35634 73724 35644 73780
rect 35700 73724 36428 73780
rect 36484 73724 42364 73780
rect 42420 73724 42430 73780
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 1362 73612 1372 73668
rect 1428 73612 7644 73668
rect 7700 73612 7710 73668
rect 8502 73612 8540 73668
rect 8596 73612 8606 73668
rect 8978 73612 8988 73668
rect 9044 73612 10332 73668
rect 10388 73612 10398 73668
rect 11330 73612 11340 73668
rect 11396 73612 15148 73668
rect 26338 73612 26348 73668
rect 26404 73612 26684 73668
rect 26740 73612 29204 73668
rect 15092 73556 15148 73612
rect 1922 73500 1932 73556
rect 1988 73500 3388 73556
rect 3444 73500 3454 73556
rect 6178 73500 6188 73556
rect 6244 73500 6972 73556
rect 7028 73500 7038 73556
rect 7858 73500 7868 73556
rect 7924 73500 14812 73556
rect 14868 73500 14878 73556
rect 15092 73500 26124 73556
rect 26180 73500 27356 73556
rect 27412 73500 28812 73556
rect 28868 73500 28878 73556
rect 29148 73444 29204 73612
rect 30482 73500 30492 73556
rect 30548 73500 37324 73556
rect 37380 73500 37390 73556
rect 6066 73388 6076 73444
rect 6132 73388 10668 73444
rect 10724 73388 10734 73444
rect 18498 73388 18508 73444
rect 18564 73388 24444 73444
rect 24500 73388 24510 73444
rect 29138 73388 29148 73444
rect 29204 73388 36876 73444
rect 36932 73388 36942 73444
rect 2034 73276 2044 73332
rect 2100 73276 5180 73332
rect 5236 73276 5246 73332
rect 6150 73276 6188 73332
rect 6244 73276 6254 73332
rect 6402 73276 6412 73332
rect 6468 73276 8316 73332
rect 8372 73276 8382 73332
rect 10210 73276 10220 73332
rect 10276 73276 11452 73332
rect 11508 73276 13020 73332
rect 13076 73276 13086 73332
rect 17686 73276 17724 73332
rect 17780 73276 17790 73332
rect 27234 73276 27244 73332
rect 27300 73276 29372 73332
rect 29428 73276 29438 73332
rect 30930 73276 30940 73332
rect 30996 73276 31500 73332
rect 31556 73276 33516 73332
rect 33572 73276 33582 73332
rect 2818 73164 2828 73220
rect 2884 73164 2940 73220
rect 2996 73164 3006 73220
rect 3714 73164 3724 73220
rect 3780 73164 4060 73220
rect 4116 73164 4126 73220
rect 4946 73164 4956 73220
rect 5012 73164 7476 73220
rect 7746 73164 7756 73220
rect 7812 73164 10108 73220
rect 10164 73164 10444 73220
rect 10500 73164 10510 73220
rect 10658 73164 10668 73220
rect 10724 73164 11788 73220
rect 11844 73164 12796 73220
rect 12852 73164 12862 73220
rect 20178 73164 20188 73220
rect 20244 73164 20860 73220
rect 20916 73164 20926 73220
rect 21074 73164 21084 73220
rect 21140 73164 22988 73220
rect 23044 73164 23054 73220
rect 25330 73164 25340 73220
rect 25396 73164 25676 73220
rect 25732 73164 25742 73220
rect 27766 73164 27804 73220
rect 27860 73164 27870 73220
rect 28802 73164 28812 73220
rect 28868 73164 29820 73220
rect 29876 73164 29886 73220
rect 32722 73164 32732 73220
rect 32788 73164 33964 73220
rect 34020 73164 34030 73220
rect 38770 73164 38780 73220
rect 38836 73164 39228 73220
rect 39284 73164 39564 73220
rect 39620 73164 39630 73220
rect 7420 73108 7476 73164
rect 4498 73052 4508 73108
rect 4564 73052 5068 73108
rect 5124 73052 5134 73108
rect 5506 73052 5516 73108
rect 5572 73052 5852 73108
rect 5908 73052 7084 73108
rect 7140 73052 7150 73108
rect 7410 73052 7420 73108
rect 7476 73052 8540 73108
rect 8596 73052 9324 73108
rect 9380 73052 12572 73108
rect 12628 73052 12638 73108
rect 17714 73052 17724 73108
rect 17780 73052 18396 73108
rect 18452 73052 18462 73108
rect 25106 73052 25116 73108
rect 25172 73052 29820 73108
rect 29876 73052 30492 73108
rect 30548 73052 30558 73108
rect 32274 73052 32284 73108
rect 32340 73052 32844 73108
rect 32900 73052 33740 73108
rect 33796 73052 35084 73108
rect 35140 73052 36316 73108
rect 36372 73052 36382 73108
rect 8418 72940 8428 72996
rect 8484 72940 8540 72996
rect 8596 72940 8606 72996
rect 11890 72940 11900 72996
rect 11956 72940 18956 72996
rect 19012 72940 19022 72996
rect 19730 72940 19740 72996
rect 19796 72940 30604 72996
rect 30660 72940 30670 72996
rect 31154 72940 31164 72996
rect 31220 72940 34748 72996
rect 34804 72940 34814 72996
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 19740 72884 19796 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 6626 72828 6636 72884
rect 6692 72828 11676 72884
rect 11732 72828 11742 72884
rect 11900 72828 19796 72884
rect 20290 72828 20300 72884
rect 20356 72828 29428 72884
rect 29698 72828 29708 72884
rect 29764 72828 30268 72884
rect 30324 72828 32900 72884
rect 35970 72828 35980 72884
rect 36036 72828 55356 72884
rect 55412 72828 55422 72884
rect 11900 72772 11956 72828
rect 29372 72772 29428 72828
rect 32844 72772 32900 72828
rect 4274 72716 4284 72772
rect 4340 72716 6076 72772
rect 6132 72716 6142 72772
rect 6290 72716 6300 72772
rect 6356 72716 8652 72772
rect 8708 72716 8718 72772
rect 8876 72716 10444 72772
rect 10500 72716 10510 72772
rect 10658 72716 10668 72772
rect 10724 72716 10892 72772
rect 10948 72716 11956 72772
rect 14242 72716 14252 72772
rect 14308 72716 19516 72772
rect 19572 72716 19582 72772
rect 24322 72716 24332 72772
rect 24388 72716 29036 72772
rect 29092 72716 29102 72772
rect 29372 72716 30940 72772
rect 30996 72716 31006 72772
rect 31826 72716 31836 72772
rect 31892 72716 32620 72772
rect 32676 72716 32686 72772
rect 32844 72716 35644 72772
rect 35700 72716 35710 72772
rect 8876 72660 8932 72716
rect 2006 72604 2044 72660
rect 2100 72604 2110 72660
rect 3714 72604 3724 72660
rect 3780 72604 6636 72660
rect 6692 72604 6702 72660
rect 7186 72604 7196 72660
rect 7252 72604 8932 72660
rect 9426 72604 9436 72660
rect 9492 72604 23772 72660
rect 23828 72604 23838 72660
rect 29782 72604 29820 72660
rect 29876 72604 29886 72660
rect 30482 72604 30492 72660
rect 30548 72604 31164 72660
rect 31220 72604 31230 72660
rect 32050 72604 32060 72660
rect 32116 72604 36428 72660
rect 36484 72604 36494 72660
rect 1474 72492 1484 72548
rect 1540 72492 3836 72548
rect 3892 72492 3902 72548
rect 5058 72492 5068 72548
rect 5124 72492 5292 72548
rect 5348 72492 5358 72548
rect 6178 72492 6188 72548
rect 6244 72492 6860 72548
rect 6916 72492 6926 72548
rect 7074 72492 7084 72548
rect 7140 72492 8204 72548
rect 8260 72492 8270 72548
rect 9090 72492 9100 72548
rect 9156 72492 11340 72548
rect 11396 72492 11406 72548
rect 12198 72492 12236 72548
rect 12292 72492 12302 72548
rect 18172 72492 18396 72548
rect 18452 72492 18462 72548
rect 23426 72492 23436 72548
rect 23492 72492 24444 72548
rect 24500 72492 28588 72548
rect 28644 72492 28812 72548
rect 28868 72492 38332 72548
rect 38388 72492 38780 72548
rect 38836 72492 38846 72548
rect 18172 72436 18228 72492
rect 3266 72380 3276 72436
rect 3332 72380 6692 72436
rect 7970 72380 7980 72436
rect 8036 72380 8540 72436
rect 8596 72380 8606 72436
rect 10210 72380 10220 72436
rect 10276 72380 11004 72436
rect 11060 72380 11070 72436
rect 12898 72380 12908 72436
rect 12964 72380 15036 72436
rect 15092 72380 15102 72436
rect 16370 72380 16380 72436
rect 16436 72380 16716 72436
rect 16772 72380 16782 72436
rect 18162 72380 18172 72436
rect 18228 72380 18238 72436
rect 18508 72380 20636 72436
rect 20692 72380 23996 72436
rect 24052 72380 24062 72436
rect 24434 72380 24444 72436
rect 24500 72380 30828 72436
rect 30884 72380 35980 72436
rect 36036 72380 36046 72436
rect 38612 72380 46620 72436
rect 46676 72380 46686 72436
rect 1932 72268 5628 72324
rect 5684 72268 5694 72324
rect 5842 72268 5852 72324
rect 5908 72268 6188 72324
rect 6244 72268 6254 72324
rect 1932 72212 1988 72268
rect 6636 72212 6692 72380
rect 18508 72324 18564 72380
rect 38612 72324 38668 72380
rect 7858 72268 7868 72324
rect 7924 72268 8204 72324
rect 8260 72268 8270 72324
rect 9986 72268 9996 72324
rect 10052 72268 10556 72324
rect 10612 72268 10622 72324
rect 11106 72268 11116 72324
rect 11172 72268 11564 72324
rect 11620 72268 11630 72324
rect 13234 72268 13244 72324
rect 13300 72268 18508 72324
rect 18564 72268 18574 72324
rect 19478 72268 19516 72324
rect 19572 72268 19582 72324
rect 20402 72268 20412 72324
rect 20468 72268 25788 72324
rect 25844 72268 25854 72324
rect 30594 72268 30604 72324
rect 30660 72268 31836 72324
rect 31892 72268 31902 72324
rect 32162 72268 32172 72324
rect 32228 72268 33852 72324
rect 33908 72268 33918 72324
rect 34738 72268 34748 72324
rect 34804 72268 35084 72324
rect 35140 72268 38668 72324
rect 1922 72156 1932 72212
rect 1988 72156 1998 72212
rect 4834 72156 4844 72212
rect 4900 72156 6300 72212
rect 6356 72156 6366 72212
rect 6636 72156 19404 72212
rect 19460 72156 19470 72212
rect 21746 72156 21756 72212
rect 21812 72156 26572 72212
rect 26628 72156 28252 72212
rect 28308 72156 30268 72212
rect 30324 72156 30334 72212
rect 36418 72156 36428 72212
rect 36484 72156 38668 72212
rect 38724 72156 38734 72212
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 5394 72044 5404 72100
rect 5460 72044 5740 72100
rect 5796 72044 5806 72100
rect 6178 72044 6188 72100
rect 6244 72044 7532 72100
rect 7588 72044 7598 72100
rect 10098 72044 10108 72100
rect 10164 72044 10668 72100
rect 10724 72044 10734 72100
rect 10882 72044 10892 72100
rect 10948 72044 12796 72100
rect 12852 72044 12862 72100
rect 36306 72044 36316 72100
rect 36372 72044 37772 72100
rect 37828 72044 37838 72100
rect 38612 72044 41356 72100
rect 41412 72044 41422 72100
rect 6188 71988 6244 72044
rect 38612 71988 38668 72044
rect 2370 71932 2380 71988
rect 2436 71932 6244 71988
rect 9762 71932 9772 71988
rect 9828 71932 13804 71988
rect 13860 71932 13870 71988
rect 16146 71932 16156 71988
rect 16212 71932 18060 71988
rect 18116 71932 18126 71988
rect 24882 71932 24892 71988
rect 24948 71932 28812 71988
rect 28868 71932 28878 71988
rect 31714 71932 31724 71988
rect 31780 71932 32396 71988
rect 32452 71932 32462 71988
rect 36866 71932 36876 71988
rect 36932 71932 38668 71988
rect 3714 71820 3724 71876
rect 3780 71820 5068 71876
rect 5124 71820 5134 71876
rect 5702 71820 5740 71876
rect 5796 71820 5806 71876
rect 5954 71820 5964 71876
rect 6020 71820 10220 71876
rect 10276 71820 10286 71876
rect 11890 71820 11900 71876
rect 11956 71820 14476 71876
rect 14532 71820 17388 71876
rect 17444 71820 17454 71876
rect 26338 71820 26348 71876
rect 26404 71820 33852 71876
rect 33908 71820 33918 71876
rect 35074 71820 35084 71876
rect 35140 71820 35532 71876
rect 35588 71820 50428 71876
rect 50484 71820 50494 71876
rect 35084 71764 35140 71820
rect 2370 71708 2380 71764
rect 2436 71708 3276 71764
rect 3332 71708 3388 71764
rect 3444 71708 3454 71764
rect 3826 71708 3836 71764
rect 3892 71708 4172 71764
rect 4228 71708 4238 71764
rect 5506 71708 5516 71764
rect 5572 71708 5964 71764
rect 6020 71708 6030 71764
rect 7186 71708 7196 71764
rect 7252 71708 7980 71764
rect 8036 71708 8046 71764
rect 9986 71708 9996 71764
rect 10052 71708 10668 71764
rect 10724 71708 11340 71764
rect 11396 71708 13468 71764
rect 13524 71708 13534 71764
rect 25666 71708 25676 71764
rect 25732 71708 27580 71764
rect 27636 71708 27646 71764
rect 29138 71708 29148 71764
rect 29204 71708 30436 71764
rect 30594 71708 30604 71764
rect 30660 71708 35140 71764
rect 37762 71708 37772 71764
rect 37828 71708 41916 71764
rect 41972 71708 41982 71764
rect 30380 71652 30436 71708
rect 1586 71596 1596 71652
rect 1652 71596 2828 71652
rect 2884 71596 2894 71652
rect 3388 71596 4732 71652
rect 4788 71596 7420 71652
rect 7476 71596 7486 71652
rect 8502 71596 8540 71652
rect 8596 71596 11676 71652
rect 11732 71596 11742 71652
rect 13346 71596 13356 71652
rect 13412 71596 14028 71652
rect 14084 71596 14094 71652
rect 18722 71596 18732 71652
rect 18788 71596 29484 71652
rect 29540 71596 29550 71652
rect 30380 71596 36876 71652
rect 36932 71596 36942 71652
rect 3388 71540 3444 71596
rect 3378 71484 3388 71540
rect 3444 71484 3454 71540
rect 4498 71484 4508 71540
rect 4564 71484 5516 71540
rect 5572 71484 5582 71540
rect 7186 71484 7196 71540
rect 7252 71484 7868 71540
rect 7924 71484 10220 71540
rect 10276 71484 10286 71540
rect 13458 71484 13468 71540
rect 13524 71484 13692 71540
rect 13748 71484 13758 71540
rect 26226 71484 26236 71540
rect 26292 71484 26572 71540
rect 26628 71484 26908 71540
rect 26964 71484 26974 71540
rect 29586 71484 29596 71540
rect 29652 71484 30044 71540
rect 30100 71484 30110 71540
rect 32918 71484 32956 71540
rect 33012 71484 33022 71540
rect 5954 71372 5964 71428
rect 6020 71372 8876 71428
rect 8932 71372 9100 71428
rect 9156 71372 9166 71428
rect 12684 71372 25340 71428
rect 25396 71372 25406 71428
rect 27010 71372 27020 71428
rect 27076 71372 29708 71428
rect 29764 71372 29774 71428
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 12684 71316 12740 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 6290 71260 6300 71316
rect 6356 71260 8092 71316
rect 8148 71260 10780 71316
rect 10836 71260 12684 71316
rect 12740 71260 12750 71316
rect 13570 71260 13580 71316
rect 13636 71260 13916 71316
rect 13972 71260 22652 71316
rect 22708 71260 22718 71316
rect 27458 71260 27468 71316
rect 27524 71260 30156 71316
rect 30212 71260 30222 71316
rect 30156 71204 30212 71260
rect 4162 71148 4172 71204
rect 4228 71148 4844 71204
rect 4900 71148 13244 71204
rect 13300 71148 13310 71204
rect 14018 71148 14028 71204
rect 14084 71148 15372 71204
rect 15428 71148 15438 71204
rect 20850 71148 20860 71204
rect 20916 71148 25228 71204
rect 25284 71148 25294 71204
rect 29558 71148 29596 71204
rect 29652 71148 29662 71204
rect 30156 71148 33404 71204
rect 33460 71148 35196 71204
rect 35252 71148 35980 71204
rect 36036 71148 36046 71204
rect 3938 71036 3948 71092
rect 4004 71036 4284 71092
rect 4340 71036 4350 71092
rect 4610 71036 4620 71092
rect 4676 71036 4956 71092
rect 5012 71036 5022 71092
rect 6402 71036 6412 71092
rect 6468 71036 8652 71092
rect 8708 71036 10892 71092
rect 10948 71036 10958 71092
rect 13794 71036 13804 71092
rect 13860 71036 23772 71092
rect 23828 71036 23838 71092
rect 29698 71036 29708 71092
rect 29764 71036 35532 71092
rect 35588 71036 35598 71092
rect 3266 70924 3276 70980
rect 3332 70924 4396 70980
rect 4452 70924 4462 70980
rect 4834 70924 4844 70980
rect 4900 70924 4956 70980
rect 5012 70924 5022 70980
rect 6290 70924 6300 70980
rect 6356 70924 6524 70980
rect 6580 70924 6590 70980
rect 7298 70924 7308 70980
rect 7364 70924 8092 70980
rect 8148 70924 12572 70980
rect 12628 70924 12638 70980
rect 13010 70924 13020 70980
rect 13076 70924 18396 70980
rect 18452 70924 18462 70980
rect 19394 70924 19404 70980
rect 19460 70924 29372 70980
rect 29428 70924 29438 70980
rect 30370 70924 30380 70980
rect 30436 70924 30884 70980
rect 31042 70924 31052 70980
rect 31108 70924 33404 70980
rect 33460 70924 33470 70980
rect 34626 70924 34636 70980
rect 34692 70924 37100 70980
rect 37156 70924 37166 70980
rect 30828 70868 30884 70924
rect 34636 70868 34692 70924
rect 2258 70812 2268 70868
rect 2324 70812 15260 70868
rect 15316 70812 15326 70868
rect 25414 70812 25452 70868
rect 25508 70812 27244 70868
rect 27300 70812 27310 70868
rect 30828 70812 34692 70868
rect 3332 70700 4956 70756
rect 5012 70700 5404 70756
rect 5460 70700 5852 70756
rect 5908 70700 5918 70756
rect 6402 70700 6412 70756
rect 6468 70700 8092 70756
rect 8148 70700 8316 70756
rect 8372 70700 8382 70756
rect 11106 70700 11116 70756
rect 11172 70700 11788 70756
rect 11844 70700 12908 70756
rect 12964 70700 12974 70756
rect 13682 70700 13692 70756
rect 13748 70700 14588 70756
rect 14644 70700 14654 70756
rect 15092 70700 17612 70756
rect 17668 70700 17678 70756
rect 20962 70700 20972 70756
rect 21028 70700 23548 70756
rect 23604 70700 23614 70756
rect 23986 70700 23996 70756
rect 24052 70700 24332 70756
rect 24388 70700 24398 70756
rect 26002 70700 26012 70756
rect 26068 70700 30380 70756
rect 30436 70700 30446 70756
rect 31714 70700 31724 70756
rect 31780 70700 32172 70756
rect 32228 70700 32238 70756
rect 33254 70700 33292 70756
rect 33348 70700 33358 70756
rect 3332 70644 3388 70700
rect 15092 70644 15148 70700
rect 1698 70588 1708 70644
rect 1764 70588 2380 70644
rect 2436 70588 3388 70644
rect 5170 70588 5180 70644
rect 5236 70588 6076 70644
rect 6132 70588 6142 70644
rect 6738 70588 6748 70644
rect 6804 70588 6860 70644
rect 6916 70588 6926 70644
rect 7410 70588 7420 70644
rect 7476 70588 8428 70644
rect 10322 70588 10332 70644
rect 10388 70588 10556 70644
rect 10612 70588 10622 70644
rect 12338 70588 12348 70644
rect 12404 70588 12460 70644
rect 12516 70588 12526 70644
rect 12674 70588 12684 70644
rect 12740 70588 14924 70644
rect 14980 70588 15148 70644
rect 15362 70588 15372 70644
rect 15428 70588 16380 70644
rect 16436 70588 16446 70644
rect 16706 70588 16716 70644
rect 16772 70588 19180 70644
rect 19236 70588 19246 70644
rect 21298 70588 21308 70644
rect 21364 70588 21644 70644
rect 21700 70588 21710 70644
rect 22866 70588 22876 70644
rect 22932 70588 23660 70644
rect 23716 70588 23726 70644
rect 23874 70588 23884 70644
rect 23940 70588 27692 70644
rect 27748 70588 37772 70644
rect 37828 70588 37838 70644
rect 8372 70532 8428 70588
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 4386 70476 4396 70532
rect 4452 70476 5964 70532
rect 6020 70476 7308 70532
rect 7364 70476 7374 70532
rect 8372 70476 16492 70532
rect 16548 70476 16558 70532
rect 16930 70476 16940 70532
rect 16996 70476 18844 70532
rect 18900 70476 18910 70532
rect 25106 70476 25116 70532
rect 25172 70476 27356 70532
rect 27412 70476 27422 70532
rect 27570 70476 27580 70532
rect 27636 70476 29372 70532
rect 29428 70476 32172 70532
rect 32228 70476 32238 70532
rect 32386 70476 32396 70532
rect 32452 70476 32462 70532
rect 32610 70476 32620 70532
rect 32676 70476 37212 70532
rect 37268 70476 37278 70532
rect 2258 70364 2268 70420
rect 2324 70364 2716 70420
rect 2772 70364 5628 70420
rect 5684 70364 5740 70420
rect 5796 70364 5806 70420
rect 6066 70364 6076 70420
rect 6132 70364 6300 70420
rect 6356 70364 6366 70420
rect 6710 70364 6748 70420
rect 6804 70364 6814 70420
rect 7522 70364 7532 70420
rect 7588 70364 8092 70420
rect 8148 70364 8316 70420
rect 8372 70364 8382 70420
rect 8530 70364 8540 70420
rect 8596 70364 8708 70420
rect 9090 70364 9100 70420
rect 9156 70364 20412 70420
rect 20468 70364 20478 70420
rect 8652 70308 8708 70364
rect 32396 70308 32452 70476
rect 32834 70364 32844 70420
rect 32900 70364 33740 70420
rect 33796 70364 33806 70420
rect 34850 70364 34860 70420
rect 34916 70364 36428 70420
rect 36484 70364 36494 70420
rect 6178 70252 6188 70308
rect 6244 70252 8428 70308
rect 8484 70252 8494 70308
rect 8652 70252 10444 70308
rect 10500 70252 10510 70308
rect 11414 70252 11452 70308
rect 11508 70252 11518 70308
rect 13682 70252 13692 70308
rect 13748 70252 18732 70308
rect 18788 70252 18798 70308
rect 24882 70252 24892 70308
rect 24948 70252 29596 70308
rect 29652 70252 29662 70308
rect 29810 70252 29820 70308
rect 29876 70252 30492 70308
rect 30548 70252 30558 70308
rect 31042 70252 31052 70308
rect 31108 70252 35084 70308
rect 35140 70252 35150 70308
rect 32284 70196 32340 70252
rect 3714 70140 3724 70196
rect 3780 70140 3836 70196
rect 3892 70140 3902 70196
rect 8194 70140 8204 70196
rect 8260 70140 9996 70196
rect 10052 70140 10062 70196
rect 11778 70140 11788 70196
rect 11844 70140 16604 70196
rect 16660 70140 16670 70196
rect 17826 70140 17836 70196
rect 17892 70140 18396 70196
rect 18452 70140 18462 70196
rect 22754 70140 22764 70196
rect 22820 70140 23212 70196
rect 23268 70140 24332 70196
rect 24388 70140 25116 70196
rect 25172 70140 25182 70196
rect 32274 70140 32284 70196
rect 32340 70140 32350 70196
rect 32498 70140 32508 70196
rect 32564 70140 35756 70196
rect 35812 70140 36988 70196
rect 37044 70140 37324 70196
rect 37380 70140 37390 70196
rect 2370 70028 2380 70084
rect 2436 70028 5180 70084
rect 5236 70028 5246 70084
rect 7270 70028 7308 70084
rect 7364 70028 7374 70084
rect 7522 70028 7532 70084
rect 7588 70028 8428 70084
rect 8484 70028 8494 70084
rect 8642 70028 8652 70084
rect 8708 70028 8764 70084
rect 8820 70028 8830 70084
rect 9426 70028 9436 70084
rect 9492 70028 13468 70084
rect 13524 70028 13534 70084
rect 17378 70028 17388 70084
rect 17444 70028 18676 70084
rect 18834 70028 18844 70084
rect 18900 70028 19516 70084
rect 19572 70028 20188 70084
rect 20244 70028 20254 70084
rect 25638 70028 25676 70084
rect 25732 70028 25742 70084
rect 26562 70028 26572 70084
rect 26628 70028 26796 70084
rect 26852 70028 26862 70084
rect 27346 70028 27356 70084
rect 27412 70028 30044 70084
rect 30100 70028 30110 70084
rect 31266 70028 31276 70084
rect 31332 70028 32060 70084
rect 32116 70028 32396 70084
rect 32452 70028 34636 70084
rect 34692 70028 35532 70084
rect 35588 70028 35598 70084
rect 18620 69972 18676 70028
rect 3042 69916 3052 69972
rect 3108 69916 5460 69972
rect 5618 69916 5628 69972
rect 5684 69916 16156 69972
rect 16212 69916 18396 69972
rect 18452 69916 18462 69972
rect 18620 69916 24892 69972
rect 24948 69916 26460 69972
rect 26516 69916 26526 69972
rect 32162 69916 32172 69972
rect 32228 69916 33516 69972
rect 33572 69916 33582 69972
rect 5404 69860 5460 69916
rect 5404 69804 9660 69860
rect 9716 69804 9726 69860
rect 9874 69804 9884 69860
rect 9940 69804 11116 69860
rect 11172 69804 11182 69860
rect 11442 69804 11452 69860
rect 11508 69804 17948 69860
rect 18004 69804 18014 69860
rect 18274 69804 18284 69860
rect 18340 69804 19628 69860
rect 19684 69804 19694 69860
rect 21298 69804 21308 69860
rect 21364 69804 27580 69860
rect 27636 69804 27646 69860
rect 30034 69804 30044 69860
rect 30100 69804 31164 69860
rect 31220 69804 32620 69860
rect 32676 69804 32686 69860
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 17948 69748 18004 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 5058 69692 5068 69748
rect 5124 69692 5628 69748
rect 5684 69692 5694 69748
rect 6626 69692 6636 69748
rect 6692 69692 9100 69748
rect 9156 69692 9166 69748
rect 9314 69692 9324 69748
rect 9380 69692 10668 69748
rect 10724 69692 10734 69748
rect 13458 69692 13468 69748
rect 13524 69692 16604 69748
rect 16660 69692 17164 69748
rect 17220 69692 17230 69748
rect 17948 69692 22540 69748
rect 22596 69692 22606 69748
rect 26002 69692 26012 69748
rect 26068 69692 35028 69748
rect 34972 69636 35028 69692
rect 3826 69580 3836 69636
rect 3892 69580 5852 69636
rect 5908 69580 5918 69636
rect 6290 69580 6300 69636
rect 6356 69580 7196 69636
rect 7252 69580 7980 69636
rect 8036 69580 8046 69636
rect 9202 69580 9212 69636
rect 9268 69580 9436 69636
rect 9492 69580 9502 69636
rect 9650 69580 9660 69636
rect 9716 69580 18172 69636
rect 18228 69580 18238 69636
rect 18470 69580 18508 69636
rect 18564 69580 18574 69636
rect 22204 69580 22988 69636
rect 23044 69580 23054 69636
rect 24322 69580 24332 69636
rect 24388 69580 28364 69636
rect 28420 69580 28430 69636
rect 28578 69580 28588 69636
rect 28644 69580 31332 69636
rect 31826 69580 31836 69636
rect 31892 69580 32732 69636
rect 32788 69580 32798 69636
rect 33506 69580 33516 69636
rect 33572 69580 34076 69636
rect 34132 69580 34142 69636
rect 34972 69580 35308 69636
rect 35364 69580 35374 69636
rect 22204 69524 22260 69580
rect 31276 69524 31332 69580
rect 1922 69468 1932 69524
rect 1988 69468 3164 69524
rect 3220 69468 4508 69524
rect 4564 69468 5404 69524
rect 5460 69468 5470 69524
rect 7420 69468 9548 69524
rect 9604 69468 12124 69524
rect 12180 69468 12190 69524
rect 12674 69468 12684 69524
rect 12740 69468 22260 69524
rect 22418 69468 22428 69524
rect 22484 69468 26180 69524
rect 26450 69468 26460 69524
rect 26516 69468 30156 69524
rect 30212 69468 31052 69524
rect 31108 69468 31118 69524
rect 31276 69468 32508 69524
rect 32564 69468 32574 69524
rect 7420 69412 7476 69468
rect 26124 69412 26180 69468
rect 3714 69356 3724 69412
rect 3780 69356 7476 69412
rect 7634 69356 7644 69412
rect 7700 69356 7868 69412
rect 7924 69356 7934 69412
rect 8194 69356 8204 69412
rect 8260 69356 9324 69412
rect 9380 69356 9390 69412
rect 9538 69356 9548 69412
rect 9604 69356 11900 69412
rect 11956 69356 13692 69412
rect 13748 69356 13758 69412
rect 18610 69356 18620 69412
rect 18676 69356 25172 69412
rect 26114 69356 26124 69412
rect 26180 69356 26190 69412
rect 27122 69356 27132 69412
rect 27188 69356 28028 69412
rect 28084 69356 28094 69412
rect 28578 69356 28588 69412
rect 28644 69356 29036 69412
rect 29092 69356 29102 69412
rect 30258 69356 30268 69412
rect 30324 69356 31724 69412
rect 31780 69356 31790 69412
rect 33394 69356 33404 69412
rect 33460 69356 34076 69412
rect 34132 69356 34142 69412
rect 9548 69300 9604 69356
rect 25116 69300 25172 69356
rect 2146 69244 2156 69300
rect 2212 69244 4284 69300
rect 4340 69244 4350 69300
rect 5702 69244 5740 69300
rect 5796 69244 5806 69300
rect 6038 69244 6076 69300
rect 6132 69244 6142 69300
rect 6626 69244 6636 69300
rect 6692 69244 9604 69300
rect 9762 69244 9772 69300
rect 9828 69244 9996 69300
rect 10052 69244 10062 69300
rect 11638 69244 11676 69300
rect 11732 69244 11742 69300
rect 16604 69244 20524 69300
rect 20580 69244 20590 69300
rect 20962 69244 20972 69300
rect 21028 69244 21308 69300
rect 21364 69244 21374 69300
rect 25106 69244 25116 69300
rect 25172 69244 28476 69300
rect 28532 69244 28542 69300
rect 30034 69244 30044 69300
rect 30100 69244 30828 69300
rect 30884 69244 30894 69300
rect 32610 69244 32620 69300
rect 32676 69244 33516 69300
rect 33572 69244 33582 69300
rect 16604 69188 16660 69244
rect 2482 69132 2492 69188
rect 2548 69132 4844 69188
rect 4900 69132 4910 69188
rect 5058 69132 5068 69188
rect 5124 69132 6524 69188
rect 6580 69132 7196 69188
rect 7252 69132 7262 69188
rect 9846 69132 9884 69188
rect 9940 69132 9950 69188
rect 10882 69132 10892 69188
rect 10948 69132 12124 69188
rect 12180 69132 12190 69188
rect 16594 69132 16604 69188
rect 16660 69132 16670 69188
rect 19292 69132 19964 69188
rect 20020 69132 20804 69188
rect 2818 69020 2828 69076
rect 2884 69020 12572 69076
rect 12628 69020 12638 69076
rect 18022 69020 18060 69076
rect 18116 69020 18126 69076
rect 19292 68964 19348 69132
rect 20748 69076 20804 69132
rect 21196 69132 22204 69188
rect 22260 69132 23100 69188
rect 23156 69132 25340 69188
rect 25396 69132 28588 69188
rect 28644 69132 28654 69188
rect 29922 69132 29932 69188
rect 29988 69132 31724 69188
rect 31780 69132 31790 69188
rect 32498 69132 32508 69188
rect 32564 69132 33964 69188
rect 34020 69132 34030 69188
rect 21196 69076 21252 69132
rect 20738 69020 20748 69076
rect 20804 69020 21196 69076
rect 21252 69020 21262 69076
rect 21746 69020 21756 69076
rect 21812 69020 26012 69076
rect 26068 69020 26078 69076
rect 28354 69020 28364 69076
rect 28420 69020 30044 69076
rect 30100 69020 31836 69076
rect 31892 69020 31902 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 4274 68908 4284 68964
rect 4340 68908 4956 68964
rect 5012 68908 5022 68964
rect 5394 68908 5404 68964
rect 5460 68908 8428 68964
rect 9426 68908 9436 68964
rect 9492 68908 10780 68964
rect 10836 68908 10846 68964
rect 12796 68908 13468 68964
rect 13524 68908 13534 68964
rect 16482 68908 16492 68964
rect 16548 68908 19292 68964
rect 19348 68908 19358 68964
rect 20178 68908 20188 68964
rect 20244 68908 26124 68964
rect 26180 68908 26572 68964
rect 26628 68908 26638 68964
rect 26786 68908 26796 68964
rect 26852 68908 26862 68964
rect 28802 68908 28812 68964
rect 28868 68908 29932 68964
rect 29988 68908 30716 68964
rect 30772 68908 30782 68964
rect 31714 68908 31724 68964
rect 31780 68908 32844 68964
rect 32900 68908 32910 68964
rect 8372 68852 8428 68908
rect 12796 68852 12852 68908
rect 26796 68852 26852 68908
rect 2370 68796 2380 68852
rect 2436 68796 3164 68852
rect 3220 68796 3230 68852
rect 3714 68796 3724 68852
rect 3780 68796 6020 68852
rect 8372 68796 8876 68852
rect 8932 68796 10108 68852
rect 10164 68796 11004 68852
rect 11060 68796 11564 68852
rect 11620 68796 12852 68852
rect 13580 68796 14980 68852
rect 15138 68796 15148 68852
rect 15204 68796 15484 68852
rect 15540 68796 15550 68852
rect 21746 68796 21756 68852
rect 21812 68796 25676 68852
rect 25732 68796 25742 68852
rect 26338 68796 26348 68852
rect 26404 68796 26852 68852
rect 28018 68796 28028 68852
rect 28084 68796 28252 68852
rect 28308 68796 28318 68852
rect 29698 68796 29708 68852
rect 29764 68796 32508 68852
rect 32564 68796 32574 68852
rect 32946 68796 32956 68852
rect 33012 68796 33852 68852
rect 33908 68796 33918 68852
rect 35522 68796 35532 68852
rect 35588 68796 40796 68852
rect 40852 68796 40862 68852
rect 5964 68740 6020 68796
rect 13580 68740 13636 68796
rect 2818 68684 2828 68740
rect 2884 68684 2940 68740
rect 2996 68684 3006 68740
rect 3378 68684 3388 68740
rect 3444 68684 3612 68740
rect 3668 68684 3678 68740
rect 3826 68684 3836 68740
rect 3892 68684 3948 68740
rect 4004 68684 4396 68740
rect 4452 68684 4462 68740
rect 5954 68684 5964 68740
rect 6020 68684 10948 68740
rect 10892 68628 10948 68684
rect 12684 68684 13636 68740
rect 14924 68740 14980 68796
rect 14924 68684 17500 68740
rect 17556 68684 17836 68740
rect 17892 68684 18172 68740
rect 18228 68684 18238 68740
rect 22092 68684 31388 68740
rect 31444 68684 31454 68740
rect 31602 68684 31612 68740
rect 31668 68684 31836 68740
rect 31892 68684 32844 68740
rect 32900 68684 32910 68740
rect 33506 68684 33516 68740
rect 33572 68684 34524 68740
rect 34580 68684 37884 68740
rect 37940 68684 37950 68740
rect 12684 68628 12740 68684
rect 2034 68572 2044 68628
rect 2100 68572 4676 68628
rect 4834 68572 4844 68628
rect 4900 68572 5068 68628
rect 5124 68572 5134 68628
rect 9650 68572 9660 68628
rect 9716 68572 10108 68628
rect 10164 68572 10174 68628
rect 10434 68572 10444 68628
rect 10500 68572 10668 68628
rect 10724 68572 10734 68628
rect 10882 68572 10892 68628
rect 10948 68572 12684 68628
rect 12740 68572 12750 68628
rect 12898 68572 12908 68628
rect 12964 68572 21868 68628
rect 21924 68572 21934 68628
rect 4620 68516 4676 68572
rect 4620 68460 6972 68516
rect 7028 68460 7038 68516
rect 8194 68460 8204 68516
rect 8260 68460 8428 68516
rect 8484 68460 8494 68516
rect 9314 68460 9324 68516
rect 9380 68460 10444 68516
rect 10500 68460 10510 68516
rect 11676 68460 21756 68516
rect 21812 68460 21822 68516
rect 1138 68348 1148 68404
rect 1204 68348 3388 68404
rect 5254 68348 5292 68404
rect 5348 68348 5358 68404
rect 7186 68348 7196 68404
rect 7252 68348 10332 68404
rect 10388 68348 10398 68404
rect 10966 68348 11004 68404
rect 11060 68348 11070 68404
rect 3332 68292 3388 68348
rect 11676 68292 11732 68460
rect 15586 68348 15596 68404
rect 15652 68348 21868 68404
rect 21924 68348 21934 68404
rect 22092 68292 22148 68684
rect 22306 68572 22316 68628
rect 22372 68572 24892 68628
rect 24948 68572 26012 68628
rect 26068 68572 26078 68628
rect 26226 68572 26236 68628
rect 26292 68572 29148 68628
rect 29204 68572 29214 68628
rect 30706 68572 30716 68628
rect 30772 68572 31500 68628
rect 31556 68572 32284 68628
rect 32340 68572 32350 68628
rect 24434 68460 24444 68516
rect 24500 68460 28700 68516
rect 28756 68460 28766 68516
rect 31378 68460 31388 68516
rect 31444 68460 32620 68516
rect 32676 68460 32686 68516
rect 34402 68460 34412 68516
rect 34468 68460 36204 68516
rect 36260 68460 36270 68516
rect 24098 68348 24108 68404
rect 24164 68348 24780 68404
rect 24836 68348 25900 68404
rect 25956 68348 25966 68404
rect 34188 68348 35308 68404
rect 35364 68348 35374 68404
rect 34188 68292 34244 68348
rect 3332 68236 4284 68292
rect 4340 68236 4350 68292
rect 4946 68236 4956 68292
rect 5012 68236 11452 68292
rect 11508 68236 11518 68292
rect 11666 68236 11676 68292
rect 11732 68236 11742 68292
rect 11890 68236 11900 68292
rect 11956 68236 16380 68292
rect 16436 68236 16446 68292
rect 16930 68236 16940 68292
rect 16996 68236 18508 68292
rect 18564 68236 22148 68292
rect 27794 68236 27804 68292
rect 27860 68236 34244 68292
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 3714 68124 3724 68180
rect 3780 68124 3836 68180
rect 3892 68124 3902 68180
rect 4834 68124 4844 68180
rect 4900 68124 9940 68180
rect 10322 68124 10332 68180
rect 10388 68124 15148 68180
rect 15204 68124 15214 68180
rect 20066 68124 20076 68180
rect 20132 68124 21196 68180
rect 21252 68124 25452 68180
rect 25508 68124 25518 68180
rect 29138 68124 29148 68180
rect 29204 68124 34188 68180
rect 34244 68124 34860 68180
rect 34916 68124 34926 68180
rect 1922 68012 1932 68068
rect 1988 68012 3164 68068
rect 3220 68012 8876 68068
rect 8932 68012 8942 68068
rect 9314 68012 9324 68068
rect 9380 68012 9436 68068
rect 9492 68012 9502 68068
rect 9884 67956 9940 68124
rect 10098 68012 10108 68068
rect 10164 68012 10444 68068
rect 10500 68012 10510 68068
rect 11732 68012 14028 68068
rect 14084 68012 17836 68068
rect 17892 68012 18284 68068
rect 18340 68012 18350 68068
rect 25554 68012 25564 68068
rect 25620 68012 29596 68068
rect 29652 68012 29662 68068
rect 11732 67956 11788 68012
rect 3378 67900 3388 67956
rect 3444 67900 9324 67956
rect 9380 67900 9390 67956
rect 9884 67900 11788 67956
rect 12674 67900 12684 67956
rect 12740 67900 15708 67956
rect 15764 67900 17164 67956
rect 17220 67900 24444 67956
rect 24500 67900 24510 67956
rect 24770 67900 24780 67956
rect 24836 67900 27356 67956
rect 27412 67900 27422 67956
rect 28802 67900 28812 67956
rect 28868 67900 29372 67956
rect 29428 67900 29820 67956
rect 29876 67900 29886 67956
rect 30594 67900 30604 67956
rect 30660 67900 31388 67956
rect 31444 67900 31454 67956
rect 2818 67788 2828 67844
rect 2884 67788 4284 67844
rect 4340 67788 4350 67844
rect 4610 67788 4620 67844
rect 4676 67788 13804 67844
rect 13860 67788 14812 67844
rect 14868 67788 14878 67844
rect 15026 67788 15036 67844
rect 15092 67788 16268 67844
rect 16324 67788 16334 67844
rect 18610 67788 18620 67844
rect 18676 67788 21420 67844
rect 21476 67788 21756 67844
rect 21812 67788 21822 67844
rect 21980 67788 22092 67844
rect 22148 67788 23436 67844
rect 23492 67788 23502 67844
rect 23874 67788 23884 67844
rect 23940 67788 24220 67844
rect 24276 67788 24286 67844
rect 27458 67788 27468 67844
rect 27524 67788 34412 67844
rect 34468 67788 34478 67844
rect 21980 67732 22036 67788
rect 3266 67676 3276 67732
rect 3332 67676 11228 67732
rect 11284 67676 11294 67732
rect 11778 67676 11788 67732
rect 11844 67676 16716 67732
rect 16772 67676 16782 67732
rect 17490 67676 17500 67732
rect 17556 67676 22036 67732
rect 22306 67676 22316 67732
rect 22372 67676 29932 67732
rect 29988 67676 33964 67732
rect 34020 67676 34030 67732
rect 11228 67620 11284 67676
rect 1922 67564 1932 67620
rect 1988 67564 3276 67620
rect 3332 67564 5068 67620
rect 5124 67564 5134 67620
rect 6514 67564 6524 67620
rect 6580 67564 7308 67620
rect 7364 67564 7374 67620
rect 11228 67564 15932 67620
rect 15988 67564 15998 67620
rect 17714 67564 17724 67620
rect 17780 67564 21980 67620
rect 22036 67564 23212 67620
rect 23268 67564 23278 67620
rect 24546 67564 24556 67620
rect 24612 67564 27580 67620
rect 27636 67564 27646 67620
rect 31938 67564 31948 67620
rect 32004 67564 32508 67620
rect 32564 67564 34412 67620
rect 34468 67564 34478 67620
rect 2034 67452 2044 67508
rect 2100 67452 5572 67508
rect 6290 67452 6300 67508
rect 6356 67452 6860 67508
rect 6916 67452 9884 67508
rect 9940 67452 9950 67508
rect 20850 67452 20860 67508
rect 20916 67452 24108 67508
rect 24164 67452 24174 67508
rect 24406 67452 24444 67508
rect 24500 67452 24510 67508
rect 25778 67452 25788 67508
rect 25844 67452 26796 67508
rect 26852 67452 26862 67508
rect 28018 67452 28028 67508
rect 28084 67452 35980 67508
rect 36036 67452 36046 67508
rect 5516 67396 5572 67452
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 2342 67340 2380 67396
rect 2436 67340 2446 67396
rect 3154 67340 3164 67396
rect 3220 67340 3276 67396
rect 3332 67340 3342 67396
rect 5516 67340 8988 67396
rect 9044 67340 9054 67396
rect 9314 67340 9324 67396
rect 9380 67340 12572 67396
rect 12628 67340 12638 67396
rect 15558 67340 15596 67396
rect 15652 67340 15662 67396
rect 21634 67340 21644 67396
rect 21700 67340 26348 67396
rect 26404 67340 26414 67396
rect 3826 67228 3836 67284
rect 3892 67228 6188 67284
rect 6244 67228 6254 67284
rect 6738 67228 6748 67284
rect 6804 67228 7868 67284
rect 7924 67228 7934 67284
rect 8866 67228 8876 67284
rect 8932 67228 9548 67284
rect 9604 67228 9614 67284
rect 10434 67228 10444 67284
rect 10500 67228 10556 67284
rect 10612 67228 10622 67284
rect 12720 67228 12796 67284
rect 12852 67228 15036 67284
rect 15092 67228 15102 67284
rect 15810 67228 15820 67284
rect 15876 67228 16828 67284
rect 16884 67228 16894 67284
rect 17490 67228 17500 67284
rect 17556 67228 17948 67284
rect 18004 67228 18014 67284
rect 18722 67228 18732 67284
rect 18788 67228 21532 67284
rect 21588 67228 21598 67284
rect 24210 67228 24220 67284
rect 24276 67228 26236 67284
rect 26292 67228 26302 67284
rect 2594 67116 2604 67172
rect 2660 67116 3164 67172
rect 3220 67116 3230 67172
rect 3714 67116 3724 67172
rect 3780 67116 4284 67172
rect 4340 67116 4350 67172
rect 4498 67116 4508 67172
rect 4564 67116 4956 67172
rect 5012 67116 5236 67172
rect 6066 67116 6076 67172
rect 6132 67116 6636 67172
rect 6692 67116 6702 67172
rect 7410 67116 7420 67172
rect 7476 67116 10668 67172
rect 10724 67116 10734 67172
rect 15148 67116 16940 67172
rect 16996 67116 17006 67172
rect 18050 67116 18060 67172
rect 18116 67116 20076 67172
rect 20132 67116 20142 67172
rect 26086 67116 26124 67172
rect 26180 67116 26190 67172
rect 27122 67116 27132 67172
rect 27188 67116 28252 67172
rect 28308 67116 28318 67172
rect 28578 67116 28588 67172
rect 28644 67116 29148 67172
rect 29204 67116 29214 67172
rect 29362 67116 29372 67172
rect 29428 67116 31388 67172
rect 31444 67116 32396 67172
rect 32452 67116 32844 67172
rect 32900 67116 32910 67172
rect 5180 67060 5236 67116
rect 15148 67060 15204 67116
rect 28588 67060 28644 67116
rect 4610 67004 4620 67060
rect 4676 67004 4956 67060
rect 5012 67004 5022 67060
rect 5180 67004 12684 67060
rect 12740 67004 12750 67060
rect 12898 67004 12908 67060
rect 12964 67004 14252 67060
rect 14308 67004 14476 67060
rect 14532 67004 14542 67060
rect 15138 67004 15148 67060
rect 15204 67004 15260 67060
rect 15316 67004 15326 67060
rect 15474 67004 15484 67060
rect 15540 67004 15596 67060
rect 15652 67004 15662 67060
rect 16566 67004 16604 67060
rect 16660 67004 16670 67060
rect 18274 67004 18284 67060
rect 18340 67004 22092 67060
rect 22148 67004 22158 67060
rect 22642 67004 22652 67060
rect 22708 67004 26796 67060
rect 26852 67004 28644 67060
rect 28802 67004 28812 67060
rect 28868 67004 29596 67060
rect 29652 67004 31276 67060
rect 31332 67004 31342 67060
rect 2930 66892 2940 66948
rect 2996 66892 3724 66948
rect 3780 66892 3790 66948
rect 4162 66892 4172 66948
rect 4228 66892 4284 66948
rect 4340 66892 4350 66948
rect 5170 66892 5180 66948
rect 5236 66892 5852 66948
rect 5908 66892 6748 66948
rect 6804 66892 6814 66948
rect 7084 66892 8988 66948
rect 9044 66892 10108 66948
rect 10164 66892 10174 66948
rect 10546 66892 10556 66948
rect 10612 66892 10668 66948
rect 10724 66892 11340 66948
rect 11396 66892 11406 66948
rect 12002 66892 12012 66948
rect 12068 66892 12236 66948
rect 12292 66892 12302 66948
rect 14242 66892 14252 66948
rect 14308 66892 14364 66948
rect 14420 66892 14430 66948
rect 16902 66892 16940 66948
rect 16996 66892 17006 66948
rect 17378 66892 17388 66948
rect 17444 66892 17836 66948
rect 17892 66892 17948 66948
rect 18004 66892 18014 66948
rect 18508 66892 20860 66948
rect 20916 66892 20926 66948
rect 23986 66892 23996 66948
rect 24052 66892 25452 66948
rect 25508 66892 25518 66948
rect 27356 66892 27916 66948
rect 27972 66892 28700 66948
rect 28756 66892 29708 66948
rect 29764 66892 33516 66948
rect 33572 66892 33582 66948
rect 7084 66836 7140 66892
rect 4284 66780 7140 66836
rect 7298 66780 7308 66836
rect 7364 66780 7644 66836
rect 7700 66780 7710 66836
rect 7858 66780 7868 66836
rect 7924 66780 8764 66836
rect 8820 66780 8830 66836
rect 9538 66780 9548 66836
rect 9604 66780 17108 66836
rect 18246 66780 18284 66836
rect 18340 66780 18350 66836
rect 4284 66500 4340 66780
rect 17052 66724 17108 66780
rect 18508 66724 18564 66892
rect 27356 66836 27412 66892
rect 27346 66780 27356 66836
rect 27412 66780 27422 66836
rect 27570 66780 27580 66836
rect 27636 66780 39116 66836
rect 39172 66780 39182 66836
rect 4946 66668 4956 66724
rect 5012 66668 9436 66724
rect 9492 66668 9502 66724
rect 9874 66668 9884 66724
rect 9940 66668 10836 66724
rect 11442 66668 11452 66724
rect 11508 66668 14028 66724
rect 14084 66668 14094 66724
rect 14364 66668 16604 66724
rect 16660 66668 16670 66724
rect 17052 66668 18564 66724
rect 18834 66668 18844 66724
rect 18900 66668 28924 66724
rect 28980 66668 28990 66724
rect 31266 66668 31276 66724
rect 31332 66668 31948 66724
rect 32004 66668 32014 66724
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 10780 66612 10836 66668
rect 14364 66612 14420 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 4946 66556 4956 66612
rect 5012 66556 5180 66612
rect 5236 66556 5964 66612
rect 6020 66556 6030 66612
rect 6412 66556 6748 66612
rect 6804 66556 7756 66612
rect 7812 66556 8372 66612
rect 8642 66556 8652 66612
rect 8708 66556 9324 66612
rect 9380 66556 10724 66612
rect 10780 66556 11116 66612
rect 11172 66556 14420 66612
rect 14578 66556 14588 66612
rect 14644 66556 17164 66612
rect 17220 66556 17230 66612
rect 18050 66556 18060 66612
rect 18116 66556 20748 66612
rect 20804 66556 22764 66612
rect 22820 66556 22830 66612
rect 24770 66556 24780 66612
rect 24836 66556 25340 66612
rect 25396 66556 26236 66612
rect 26292 66556 26302 66612
rect 6412 66500 6468 66556
rect 8316 66500 8372 66556
rect 2706 66444 2716 66500
rect 2772 66444 2940 66500
rect 2996 66444 3006 66500
rect 3154 66444 3164 66500
rect 3220 66444 4340 66500
rect 4498 66444 4508 66500
rect 4564 66444 6468 66500
rect 6626 66444 6636 66500
rect 6692 66444 8092 66500
rect 8148 66444 8158 66500
rect 8306 66444 8316 66500
rect 8372 66444 8382 66500
rect 10668 66388 10724 66556
rect 10882 66444 10892 66500
rect 10948 66444 18732 66500
rect 18788 66444 18798 66500
rect 19954 66444 19964 66500
rect 20020 66444 21868 66500
rect 21924 66444 23548 66500
rect 23604 66444 23614 66500
rect 26114 66444 26124 66500
rect 26180 66444 35532 66500
rect 35588 66444 35598 66500
rect 2594 66332 2604 66388
rect 2660 66332 3388 66388
rect 4050 66332 4060 66388
rect 4116 66332 7868 66388
rect 7924 66332 10612 66388
rect 10668 66332 11116 66388
rect 11172 66332 11182 66388
rect 13654 66332 13692 66388
rect 13748 66332 13758 66388
rect 15026 66332 15036 66388
rect 15092 66332 19292 66388
rect 19348 66332 19358 66388
rect 20066 66332 20076 66388
rect 20132 66332 22092 66388
rect 22148 66332 22158 66388
rect 22642 66332 22652 66388
rect 22708 66332 27020 66388
rect 27076 66332 27086 66388
rect 28354 66332 28364 66388
rect 28420 66332 40348 66388
rect 40404 66332 40414 66388
rect 3332 66276 3388 66332
rect 10556 66276 10612 66332
rect 3332 66220 6636 66276
rect 6692 66220 6702 66276
rect 7158 66220 7196 66276
rect 7252 66220 7262 66276
rect 9062 66220 9100 66276
rect 9156 66220 9166 66276
rect 10546 66220 10556 66276
rect 10612 66220 15708 66276
rect 15764 66220 15774 66276
rect 15932 66220 18620 66276
rect 18676 66220 18686 66276
rect 19170 66220 19180 66276
rect 19236 66220 20300 66276
rect 20356 66220 22596 66276
rect 25442 66220 25452 66276
rect 25508 66220 26908 66276
rect 26964 66220 26974 66276
rect 27122 66220 27132 66276
rect 27188 66220 29596 66276
rect 29652 66220 29662 66276
rect 15932 66164 15988 66220
rect 22540 66164 22596 66220
rect 4274 66108 4284 66164
rect 4340 66108 6860 66164
rect 6916 66108 8876 66164
rect 8932 66108 8942 66164
rect 9426 66108 9436 66164
rect 9492 66108 11284 66164
rect 11554 66108 11564 66164
rect 11620 66108 11676 66164
rect 11732 66108 11742 66164
rect 14354 66108 14364 66164
rect 14420 66108 14812 66164
rect 14868 66108 15988 66164
rect 17826 66108 17836 66164
rect 17892 66108 22316 66164
rect 22372 66108 22382 66164
rect 22540 66108 25564 66164
rect 25620 66108 25630 66164
rect 11228 66052 11284 66108
rect 4386 65996 4396 66052
rect 4452 65996 6636 66052
rect 6692 65996 6702 66052
rect 7074 65996 7084 66052
rect 7140 65996 7532 66052
rect 7588 65996 9660 66052
rect 9716 65996 9726 66052
rect 11228 65996 12796 66052
rect 12852 65996 12862 66052
rect 14018 65996 14028 66052
rect 14084 65996 16044 66052
rect 16100 65996 16110 66052
rect 17938 65996 17948 66052
rect 18004 65996 20300 66052
rect 20356 65996 20366 66052
rect 20626 65996 20636 66052
rect 20692 65996 21756 66052
rect 21812 65996 22204 66052
rect 22260 65996 22270 66052
rect 22754 65996 22764 66052
rect 22820 65996 23436 66052
rect 23492 65996 23502 66052
rect 26002 65996 26012 66052
rect 26068 65996 27804 66052
rect 27860 65996 27870 66052
rect 1922 65884 1932 65940
rect 1988 65884 3612 65940
rect 3668 65884 4620 65940
rect 4676 65884 4686 65940
rect 4946 65884 4956 65940
rect 5012 65884 8316 65940
rect 8372 65884 8382 65940
rect 8754 65884 8764 65940
rect 8820 65884 10556 65940
rect 10612 65884 11676 65940
rect 11732 65884 15260 65940
rect 15316 65884 15326 65940
rect 21858 65884 21868 65940
rect 21924 65884 22540 65940
rect 22596 65884 24892 65940
rect 24948 65884 24958 65940
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 3714 65772 3724 65828
rect 3780 65772 4508 65828
rect 4564 65772 4574 65828
rect 5058 65772 5068 65828
rect 5124 65772 5516 65828
rect 5572 65772 15820 65828
rect 15876 65772 15886 65828
rect 20178 65772 20188 65828
rect 20244 65772 29372 65828
rect 29428 65772 29438 65828
rect 29922 65772 29932 65828
rect 29988 65772 30604 65828
rect 30660 65772 30670 65828
rect 3042 65660 3052 65716
rect 3108 65660 5628 65716
rect 5684 65660 5694 65716
rect 5842 65660 5852 65716
rect 5908 65660 6076 65716
rect 6132 65660 6524 65716
rect 6580 65660 6590 65716
rect 7186 65660 7196 65716
rect 7252 65660 7644 65716
rect 7700 65660 7710 65716
rect 7970 65660 7980 65716
rect 8036 65660 8092 65716
rect 8148 65660 8158 65716
rect 8278 65660 8316 65716
rect 8372 65660 8382 65716
rect 12422 65660 12460 65716
rect 12516 65660 12526 65716
rect 17490 65660 17500 65716
rect 17556 65660 17948 65716
rect 18004 65660 18014 65716
rect 18134 65660 18172 65716
rect 18228 65660 18238 65716
rect 19618 65660 19628 65716
rect 19684 65660 20860 65716
rect 20916 65660 20926 65716
rect 25106 65660 25116 65716
rect 25172 65660 25452 65716
rect 25508 65660 26684 65716
rect 26740 65660 26750 65716
rect 26852 65660 27356 65716
rect 27412 65660 27422 65716
rect 28018 65660 28028 65716
rect 28084 65660 28588 65716
rect 28644 65660 29708 65716
rect 29764 65660 30492 65716
rect 30548 65660 31052 65716
rect 31108 65660 31118 65716
rect 26852 65604 26908 65660
rect 1922 65548 1932 65604
rect 1988 65548 4844 65604
rect 4900 65548 4910 65604
rect 5394 65548 5404 65604
rect 5460 65548 8204 65604
rect 8260 65548 8270 65604
rect 10434 65548 10444 65604
rect 10500 65548 16268 65604
rect 16324 65548 16334 65604
rect 20962 65548 20972 65604
rect 21028 65548 21868 65604
rect 21924 65548 21934 65604
rect 22502 65548 22540 65604
rect 22596 65548 22606 65604
rect 24882 65548 24892 65604
rect 24948 65548 26908 65604
rect 27244 65548 27468 65604
rect 27524 65548 27534 65604
rect 30370 65548 30380 65604
rect 30436 65548 31276 65604
rect 31332 65548 31342 65604
rect 2258 65436 2268 65492
rect 2324 65436 3836 65492
rect 3892 65436 3902 65492
rect 4050 65436 4060 65492
rect 4116 65436 8764 65492
rect 8820 65436 8830 65492
rect 11218 65436 11228 65492
rect 11284 65436 11452 65492
rect 11508 65436 11518 65492
rect 13010 65436 13020 65492
rect 13076 65436 14812 65492
rect 14868 65436 14878 65492
rect 15586 65436 15596 65492
rect 15652 65436 16604 65492
rect 16660 65436 16670 65492
rect 16818 65436 16828 65492
rect 16884 65436 19068 65492
rect 19124 65436 19134 65492
rect 24210 65436 24220 65492
rect 24276 65436 26012 65492
rect 26068 65436 26078 65492
rect 26450 65436 26460 65492
rect 26516 65436 27020 65492
rect 27076 65436 27086 65492
rect 26012 65380 26068 65436
rect 27244 65380 27300 65548
rect 27570 65436 27580 65492
rect 27636 65436 28140 65492
rect 28196 65436 30268 65492
rect 30324 65436 30334 65492
rect 3042 65324 3052 65380
rect 3108 65324 5740 65380
rect 5796 65324 5806 65380
rect 6626 65324 6636 65380
rect 6692 65324 9436 65380
rect 9492 65324 9502 65380
rect 10210 65324 10220 65380
rect 10276 65324 11900 65380
rect 11956 65324 13804 65380
rect 13860 65324 13916 65380
rect 13972 65324 13982 65380
rect 15092 65324 15596 65380
rect 15652 65324 15662 65380
rect 16258 65324 16268 65380
rect 16324 65324 16492 65380
rect 16548 65324 20188 65380
rect 20244 65324 20254 65380
rect 23762 65324 23772 65380
rect 23828 65324 24892 65380
rect 24948 65324 24958 65380
rect 26012 65324 26348 65380
rect 26404 65324 26414 65380
rect 26674 65324 26684 65380
rect 26740 65324 27300 65380
rect 28914 65324 28924 65380
rect 28980 65324 29484 65380
rect 29540 65324 31500 65380
rect 31556 65324 31566 65380
rect 15092 65268 15148 65324
rect 3826 65212 3836 65268
rect 3892 65212 4844 65268
rect 4900 65212 4910 65268
rect 5506 65212 5516 65268
rect 5572 65212 10108 65268
rect 10164 65212 10174 65268
rect 10322 65212 10332 65268
rect 10388 65212 15148 65268
rect 16258 65212 16268 65268
rect 16324 65212 16716 65268
rect 16772 65212 18508 65268
rect 18564 65212 18574 65268
rect 20514 65212 20524 65268
rect 20580 65212 24444 65268
rect 24500 65212 24510 65268
rect 2706 65100 2716 65156
rect 2772 65100 3052 65156
rect 3108 65100 3724 65156
rect 3780 65100 3790 65156
rect 6412 65100 6748 65156
rect 6804 65100 8540 65156
rect 8596 65100 8606 65156
rect 8754 65100 8764 65156
rect 8820 65100 19180 65156
rect 19236 65100 19246 65156
rect 23660 65100 25116 65156
rect 25172 65100 25182 65156
rect 26338 65100 26348 65156
rect 26404 65100 28812 65156
rect 28868 65100 28878 65156
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 6412 65044 6468 65100
rect 23660 65044 23716 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 4946 64988 4956 65044
rect 5012 64988 6468 65044
rect 6626 64988 6636 65044
rect 6692 64988 10108 65044
rect 10164 64988 10332 65044
rect 10388 64988 10398 65044
rect 15922 64988 15932 65044
rect 15988 64988 16492 65044
rect 16548 64988 16558 65044
rect 18386 64988 18396 65044
rect 18452 64988 23716 65044
rect 23874 64988 23884 65044
rect 23940 64988 26908 65044
rect 26964 64988 27468 65044
rect 27524 64988 27534 65044
rect 3154 64876 3164 64932
rect 3220 64876 8204 64932
rect 8260 64876 8270 64932
rect 8530 64876 8540 64932
rect 8596 64876 12460 64932
rect 12516 64876 12526 64932
rect 12898 64876 12908 64932
rect 12964 64876 13580 64932
rect 13636 64876 13646 64932
rect 14018 64876 14028 64932
rect 14084 64876 14252 64932
rect 14308 64876 14318 64932
rect 15362 64876 15372 64932
rect 15428 64876 17500 64932
rect 17556 64876 17566 64932
rect 21522 64876 21532 64932
rect 21588 64876 23548 64932
rect 23604 64876 23772 64932
rect 23828 64876 25900 64932
rect 25956 64876 25966 64932
rect 27010 64876 27020 64932
rect 27076 64876 28364 64932
rect 28420 64876 28430 64932
rect 2370 64764 2380 64820
rect 2436 64764 2828 64820
rect 2884 64764 2894 64820
rect 4946 64764 4956 64820
rect 5012 64764 5964 64820
rect 6020 64764 6030 64820
rect 6290 64764 6300 64820
rect 6356 64764 8540 64820
rect 8596 64764 10220 64820
rect 10276 64764 10444 64820
rect 10500 64764 13468 64820
rect 13524 64764 15484 64820
rect 15540 64764 15550 64820
rect 15810 64764 15820 64820
rect 15876 64764 18284 64820
rect 18340 64764 18350 64820
rect 19730 64764 19740 64820
rect 19796 64764 20524 64820
rect 20580 64764 20590 64820
rect 22418 64764 22428 64820
rect 22484 64764 23100 64820
rect 23156 64764 23324 64820
rect 23380 64764 23390 64820
rect 23986 64764 23996 64820
rect 24052 64764 25676 64820
rect 25732 64764 25742 64820
rect 28242 64764 28252 64820
rect 28308 64764 29820 64820
rect 29876 64764 29886 64820
rect 2258 64652 2268 64708
rect 2324 64652 3164 64708
rect 3220 64652 3276 64708
rect 3332 64652 3342 64708
rect 3602 64652 3612 64708
rect 3668 64652 7196 64708
rect 7252 64652 7262 64708
rect 8978 64652 8988 64708
rect 9044 64652 12124 64708
rect 12180 64652 12908 64708
rect 12964 64652 12974 64708
rect 13906 64652 13916 64708
rect 13972 64652 15036 64708
rect 15092 64652 15102 64708
rect 15922 64652 15932 64708
rect 15988 64652 17164 64708
rect 17220 64652 18508 64708
rect 18564 64652 18574 64708
rect 18722 64652 18732 64708
rect 18788 64652 23884 64708
rect 23940 64652 23950 64708
rect 25106 64652 25116 64708
rect 25172 64652 26684 64708
rect 26740 64652 26750 64708
rect 2818 64540 2828 64596
rect 2884 64540 3052 64596
rect 3108 64540 3118 64596
rect 4498 64540 4508 64596
rect 4564 64540 4956 64596
rect 5012 64540 5022 64596
rect 5170 64540 5180 64596
rect 5236 64540 6300 64596
rect 6356 64540 6366 64596
rect 7634 64540 7644 64596
rect 7700 64540 10108 64596
rect 10164 64540 10174 64596
rect 12338 64540 12348 64596
rect 12404 64540 15148 64596
rect 16370 64540 16380 64596
rect 16436 64540 18396 64596
rect 18452 64540 18462 64596
rect 21186 64540 21196 64596
rect 21252 64540 22092 64596
rect 22148 64540 22158 64596
rect 25442 64540 25452 64596
rect 25508 64540 25676 64596
rect 25732 64540 25742 64596
rect 3378 64428 3388 64484
rect 3444 64428 4060 64484
rect 4116 64428 4126 64484
rect 4834 64428 4844 64484
rect 4900 64428 7476 64484
rect 7830 64428 7868 64484
rect 7924 64428 7934 64484
rect 8978 64428 8988 64484
rect 9044 64428 12236 64484
rect 12292 64428 12302 64484
rect 12562 64428 12572 64484
rect 12628 64428 13916 64484
rect 13972 64428 13982 64484
rect 7420 64372 7476 64428
rect 15092 64372 15148 64540
rect 17164 64484 17220 64540
rect 16034 64428 16044 64484
rect 16100 64428 16604 64484
rect 16660 64428 16670 64484
rect 17154 64428 17164 64484
rect 17220 64428 17230 64484
rect 17602 64428 17612 64484
rect 17668 64428 19852 64484
rect 19908 64428 19918 64484
rect 22418 64428 22428 64484
rect 22484 64428 24332 64484
rect 24388 64428 24398 64484
rect 6962 64316 6972 64372
rect 7028 64316 7196 64372
rect 7252 64316 7262 64372
rect 7420 64316 8092 64372
rect 8148 64316 8158 64372
rect 8754 64316 8764 64372
rect 8820 64316 10444 64372
rect 10500 64316 10510 64372
rect 15092 64316 18172 64372
rect 18228 64316 18732 64372
rect 18788 64316 18798 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 2370 64204 2380 64260
rect 2436 64204 11452 64260
rect 11508 64204 13580 64260
rect 13636 64204 15260 64260
rect 15316 64204 15326 64260
rect 15474 64204 15484 64260
rect 15540 64204 19628 64260
rect 19684 64204 19694 64260
rect 22978 64204 22988 64260
rect 23044 64204 23436 64260
rect 23492 64204 23502 64260
rect 24882 64204 24892 64260
rect 24948 64204 26684 64260
rect 26740 64204 26750 64260
rect 2146 64092 2156 64148
rect 2212 64092 4956 64148
rect 5012 64092 5022 64148
rect 5506 64092 5516 64148
rect 5572 64092 9100 64148
rect 9156 64092 9166 64148
rect 12226 64092 12236 64148
rect 12292 64092 13132 64148
rect 13188 64092 13692 64148
rect 13748 64092 13758 64148
rect 13990 64092 14028 64148
rect 14084 64092 14094 64148
rect 15138 64092 15148 64148
rect 15204 64092 16828 64148
rect 16884 64092 18284 64148
rect 18340 64092 18350 64148
rect 18946 64092 18956 64148
rect 19012 64092 19740 64148
rect 19796 64092 20300 64148
rect 20356 64092 20366 64148
rect 20850 64092 20860 64148
rect 20916 64092 22204 64148
rect 22260 64092 24108 64148
rect 24164 64092 24174 64148
rect 26562 64092 26572 64148
rect 26628 64092 27132 64148
rect 27188 64092 28924 64148
rect 28980 64092 28990 64148
rect 13692 64036 13748 64092
rect 1810 63980 1820 64036
rect 1876 63980 3612 64036
rect 3668 63980 3678 64036
rect 3826 63980 3836 64036
rect 3892 63980 3948 64036
rect 4004 63980 4014 64036
rect 4956 63980 8652 64036
rect 8708 63980 8718 64036
rect 11900 63980 12908 64036
rect 12964 63980 12974 64036
rect 13692 63980 15708 64036
rect 15764 63980 15774 64036
rect 17042 63980 17052 64036
rect 17108 63980 17118 64036
rect 18834 63980 18844 64036
rect 18900 63980 20188 64036
rect 20244 63980 20254 64036
rect 21298 63980 21308 64036
rect 21364 63980 21374 64036
rect 23426 63980 23436 64036
rect 23492 63980 25788 64036
rect 25844 63980 28252 64036
rect 28308 63980 28318 64036
rect 4956 63924 5012 63980
rect 11900 63924 11956 63980
rect 17052 63924 17108 63980
rect 21308 63924 21364 63980
rect 27132 63924 27188 63980
rect 2370 63868 2380 63924
rect 2436 63868 3276 63924
rect 3332 63868 3342 63924
rect 3714 63868 3724 63924
rect 3780 63868 5012 63924
rect 6850 63868 6860 63924
rect 6916 63868 9996 63924
rect 10052 63868 10062 63924
rect 10332 63868 11228 63924
rect 11284 63868 11294 63924
rect 11890 63868 11900 63924
rect 11956 63868 11966 63924
rect 12562 63868 12572 63924
rect 12628 63868 15484 63924
rect 15540 63868 15550 63924
rect 17052 63868 18172 63924
rect 18228 63868 18238 63924
rect 18320 63868 18396 63924
rect 18452 63868 18462 63924
rect 18722 63868 18732 63924
rect 18788 63868 19292 63924
rect 19348 63868 19358 63924
rect 19618 63868 19628 63924
rect 19684 63868 20300 63924
rect 20356 63868 21364 63924
rect 22194 63868 22204 63924
rect 22260 63868 22988 63924
rect 23044 63868 23054 63924
rect 23874 63868 23884 63924
rect 23940 63868 26460 63924
rect 26516 63868 26526 63924
rect 26674 63868 26684 63924
rect 26740 63868 26908 63924
rect 26964 63868 26974 63924
rect 27122 63868 27132 63924
rect 27188 63868 27198 63924
rect 10332 63812 10388 63868
rect 18396 63812 18452 63868
rect 1922 63756 1932 63812
rect 1988 63756 3164 63812
rect 3220 63756 4844 63812
rect 4900 63756 4910 63812
rect 6290 63756 6300 63812
rect 6356 63756 7084 63812
rect 7140 63756 7980 63812
rect 8036 63756 8046 63812
rect 8418 63756 8428 63812
rect 8484 63756 10220 63812
rect 10276 63756 10332 63812
rect 10388 63756 10398 63812
rect 11330 63756 11340 63812
rect 11396 63756 12348 63812
rect 12404 63756 12414 63812
rect 17042 63756 17052 63812
rect 17108 63756 17612 63812
rect 17668 63756 17724 63812
rect 17780 63756 17790 63812
rect 18396 63756 19180 63812
rect 19236 63756 19246 63812
rect 25890 63756 25900 63812
rect 25956 63756 26684 63812
rect 26740 63756 26750 63812
rect 26898 63756 26908 63812
rect 26964 63756 38332 63812
rect 38388 63756 38398 63812
rect 2370 63644 2380 63700
rect 2436 63644 3388 63700
rect 4162 63644 4172 63700
rect 4228 63644 7756 63700
rect 7812 63644 8540 63700
rect 8596 63644 8606 63700
rect 9202 63644 9212 63700
rect 9268 63644 9548 63700
rect 9604 63644 16604 63700
rect 16660 63644 17388 63700
rect 17444 63644 17454 63700
rect 18610 63644 18620 63700
rect 18676 63644 18956 63700
rect 19012 63644 20636 63700
rect 20692 63644 21308 63700
rect 21364 63644 23660 63700
rect 23716 63644 23726 63700
rect 24210 63644 24220 63700
rect 24276 63644 25116 63700
rect 25172 63644 25182 63700
rect 2482 63532 2492 63588
rect 2548 63532 3164 63588
rect 3220 63532 3230 63588
rect 3332 63476 3388 63644
rect 7232 63532 7308 63588
rect 7364 63532 7644 63588
rect 7700 63532 8764 63588
rect 8820 63532 11788 63588
rect 11844 63532 12012 63588
rect 12068 63532 12078 63588
rect 22306 63532 22316 63588
rect 22372 63532 23324 63588
rect 23380 63532 24780 63588
rect 24836 63532 24846 63588
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 2678 63420 2716 63476
rect 2772 63420 2782 63476
rect 3332 63420 3500 63476
rect 3556 63420 3566 63476
rect 7186 63420 7196 63476
rect 7252 63420 8204 63476
rect 8260 63420 9268 63476
rect 9986 63420 9996 63476
rect 10052 63420 15148 63476
rect 15250 63420 15260 63476
rect 15316 63420 16044 63476
rect 16100 63420 16110 63476
rect 16268 63420 23212 63476
rect 23268 63420 23278 63476
rect 24098 63420 24108 63476
rect 24164 63420 24556 63476
rect 24612 63420 24622 63476
rect 9212 63364 9268 63420
rect 15092 63364 15148 63420
rect 16268 63364 16324 63420
rect 3574 63308 3612 63364
rect 3668 63308 3678 63364
rect 4162 63308 4172 63364
rect 4228 63308 7308 63364
rect 7364 63308 7374 63364
rect 7532 63308 7980 63364
rect 8036 63308 8876 63364
rect 8932 63308 8942 63364
rect 9212 63308 11340 63364
rect 11396 63308 11406 63364
rect 11526 63308 11564 63364
rect 11620 63308 11630 63364
rect 15092 63308 16324 63364
rect 16640 63308 16716 63364
rect 16772 63308 18620 63364
rect 18676 63308 18686 63364
rect 21970 63308 21980 63364
rect 22036 63308 22876 63364
rect 22932 63308 23884 63364
rect 23940 63308 23950 63364
rect 24322 63308 24332 63364
rect 24388 63308 25172 63364
rect 7532 63252 7588 63308
rect 4610 63196 4620 63252
rect 4676 63196 5852 63252
rect 5908 63196 6636 63252
rect 6692 63196 6702 63252
rect 6850 63196 6860 63252
rect 6916 63196 7588 63252
rect 8306 63196 8316 63252
rect 8372 63196 9996 63252
rect 10052 63196 10062 63252
rect 14018 63196 14028 63252
rect 14084 63196 15260 63252
rect 15316 63196 15326 63252
rect 15698 63196 15708 63252
rect 15764 63196 16380 63252
rect 16436 63196 16446 63252
rect 20402 63196 20412 63252
rect 20468 63196 21756 63252
rect 21812 63196 21822 63252
rect 23650 63196 23660 63252
rect 23716 63196 24220 63252
rect 24276 63196 24286 63252
rect 25116 63140 25172 63308
rect 26852 63196 34300 63252
rect 34356 63196 34366 63252
rect 2370 63084 2380 63140
rect 2436 63084 6188 63140
rect 6244 63084 6254 63140
rect 7858 63084 7868 63140
rect 7924 63084 9212 63140
rect 9268 63084 9278 63140
rect 10098 63084 10108 63140
rect 10164 63084 10780 63140
rect 10836 63084 11788 63140
rect 12226 63084 12236 63140
rect 12292 63084 14364 63140
rect 14420 63084 15596 63140
rect 15652 63084 15662 63140
rect 21858 63084 21868 63140
rect 21924 63084 22764 63140
rect 22820 63084 22830 63140
rect 25106 63084 25116 63140
rect 25172 63084 25182 63140
rect 11732 63028 11788 63084
rect 26852 63028 26908 63196
rect 27570 63084 27580 63140
rect 27636 63084 28252 63140
rect 28308 63084 28812 63140
rect 28868 63084 29932 63140
rect 29988 63084 29998 63140
rect 4274 62972 4284 63028
rect 4340 62972 8820 63028
rect 8978 62972 8988 63028
rect 9044 62972 10556 63028
rect 10612 62972 10622 63028
rect 11732 62972 13412 63028
rect 13570 62972 13580 63028
rect 13636 62972 13692 63028
rect 13748 62972 13758 63028
rect 15250 62972 15260 63028
rect 15316 62972 16716 63028
rect 16772 62972 19740 63028
rect 19796 62972 26908 63028
rect 28466 62972 28476 63028
rect 28532 62972 29596 63028
rect 29652 62972 29662 63028
rect 8764 62916 8820 62972
rect 13356 62916 13412 62972
rect 3332 62860 6300 62916
rect 6356 62860 6366 62916
rect 7298 62860 7308 62916
rect 7364 62860 7756 62916
rect 7812 62860 8428 62916
rect 8484 62860 8494 62916
rect 8764 62860 9324 62916
rect 9380 62860 12124 62916
rect 12180 62860 12796 62916
rect 12852 62860 12862 62916
rect 13356 62860 13748 62916
rect 3332 62804 3388 62860
rect 13692 62804 13748 62860
rect 2706 62748 2716 62804
rect 2772 62748 2884 62804
rect 3154 62748 3164 62804
rect 3220 62748 3388 62804
rect 4498 62748 4508 62804
rect 4564 62748 11116 62804
rect 11172 62748 11564 62804
rect 11620 62748 13356 62804
rect 13412 62748 13422 62804
rect 13682 62748 13692 62804
rect 13748 62748 13758 62804
rect 2594 62636 2604 62692
rect 2660 62636 2670 62692
rect 2604 62244 2660 62636
rect 2828 62356 2884 62748
rect 3266 62636 3276 62692
rect 3332 62636 4844 62692
rect 4900 62636 4910 62692
rect 8530 62636 8540 62692
rect 8596 62636 10220 62692
rect 10276 62636 10286 62692
rect 11862 62636 11900 62692
rect 11956 62636 11966 62692
rect 13010 62636 13020 62692
rect 13076 62636 15596 62692
rect 15652 62636 15662 62692
rect 15810 62636 15820 62692
rect 15876 62636 17948 62692
rect 18004 62636 18014 62692
rect 19628 62580 19684 62972
rect 20850 62860 20860 62916
rect 20916 62860 21532 62916
rect 21588 62860 21598 62916
rect 21746 62860 21756 62916
rect 21812 62860 23212 62916
rect 23268 62860 26796 62916
rect 26852 62860 27692 62916
rect 27748 62860 30380 62916
rect 30436 62860 30446 62916
rect 21074 62748 21084 62804
rect 21140 62748 22092 62804
rect 22148 62748 22540 62804
rect 22596 62748 22606 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 20850 62636 20860 62692
rect 20916 62636 23660 62692
rect 23716 62636 24220 62692
rect 24276 62636 24668 62692
rect 24724 62636 25900 62692
rect 25956 62636 26348 62692
rect 26404 62636 26414 62692
rect 3332 62524 6244 62580
rect 6402 62524 6412 62580
rect 6468 62524 7420 62580
rect 7476 62524 7644 62580
rect 7700 62524 7710 62580
rect 8082 62524 8092 62580
rect 8148 62524 10780 62580
rect 10836 62524 10846 62580
rect 15250 62524 15260 62580
rect 15316 62524 16716 62580
rect 16772 62524 17612 62580
rect 17668 62524 17678 62580
rect 19628 62524 19740 62580
rect 19796 62524 19806 62580
rect 21494 62524 21532 62580
rect 21588 62524 22092 62580
rect 22148 62524 22158 62580
rect 28354 62524 28364 62580
rect 28420 62524 28812 62580
rect 28868 62524 28878 62580
rect 3332 62468 3388 62524
rect 3154 62412 3164 62468
rect 3220 62412 3388 62468
rect 6188 62468 6244 62524
rect 6188 62412 10668 62468
rect 10724 62412 10734 62468
rect 11004 62412 12236 62468
rect 12292 62412 12302 62468
rect 13346 62412 13356 62468
rect 13412 62412 15148 62468
rect 17154 62412 17164 62468
rect 17220 62412 17276 62468
rect 17332 62412 17342 62468
rect 21970 62412 21980 62468
rect 22036 62412 22204 62468
rect 22260 62412 22270 62468
rect 11004 62356 11060 62412
rect 15092 62356 15148 62412
rect 2818 62300 2828 62356
rect 2884 62300 2894 62356
rect 3042 62300 3052 62356
rect 3108 62300 4956 62356
rect 5012 62300 5292 62356
rect 5348 62300 5358 62356
rect 5740 62300 11060 62356
rect 11218 62300 11228 62356
rect 11284 62300 13580 62356
rect 13636 62300 13646 62356
rect 15092 62300 18172 62356
rect 18228 62300 18238 62356
rect 19506 62300 19516 62356
rect 19572 62300 20860 62356
rect 20916 62300 20926 62356
rect 5740 62244 5796 62300
rect 2594 62188 2604 62244
rect 2660 62188 2670 62244
rect 2828 62188 3388 62244
rect 3444 62188 3454 62244
rect 3938 62188 3948 62244
rect 4004 62188 4172 62244
rect 4228 62188 5796 62244
rect 8194 62188 8204 62244
rect 8260 62188 8876 62244
rect 8932 62188 8942 62244
rect 9202 62188 9212 62244
rect 9268 62188 9996 62244
rect 10052 62188 10062 62244
rect 10658 62188 10668 62244
rect 10724 62188 14028 62244
rect 14084 62188 14094 62244
rect 17164 62188 19292 62244
rect 19348 62188 19628 62244
rect 19684 62188 19694 62244
rect 20132 62188 21980 62244
rect 22036 62188 22046 62244
rect 22642 62188 22652 62244
rect 22708 62188 24780 62244
rect 24836 62188 25340 62244
rect 25396 62188 25406 62244
rect 2818 62132 2828 62188
rect 2884 62132 2894 62188
rect 17164 62132 17220 62188
rect 20132 62132 20188 62188
rect 4834 62076 4844 62132
rect 4900 62076 5068 62132
rect 5124 62076 5134 62132
rect 6066 62076 6076 62132
rect 6132 62076 9772 62132
rect 9828 62076 9996 62132
rect 10052 62076 10062 62132
rect 10770 62076 10780 62132
rect 10836 62076 12012 62132
rect 12068 62076 12078 62132
rect 14354 62076 14364 62132
rect 14420 62076 15708 62132
rect 15764 62076 15774 62132
rect 16034 62076 16044 62132
rect 16100 62076 17164 62132
rect 17220 62076 17230 62132
rect 18834 62076 18844 62132
rect 18900 62076 20188 62132
rect 23548 62020 23604 62188
rect 9538 61964 9548 62020
rect 9604 61964 12908 62020
rect 12964 61964 13692 62020
rect 13748 61964 13758 62020
rect 15922 61964 15932 62020
rect 15988 61964 16380 62020
rect 16436 61964 16446 62020
rect 16818 61964 16828 62020
rect 16884 61964 17500 62020
rect 17556 61964 17566 62020
rect 18694 61964 18732 62020
rect 18788 61964 18798 62020
rect 23538 61964 23548 62020
rect 23604 61964 23614 62020
rect 23762 61964 23772 62020
rect 23828 61964 24892 62020
rect 24948 61964 24958 62020
rect 25106 61964 25116 62020
rect 25172 61964 33292 62020
rect 33348 61964 33358 62020
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 6850 61852 6860 61908
rect 6916 61852 7532 61908
rect 7588 61852 7598 61908
rect 10546 61852 10556 61908
rect 10612 61852 13804 61908
rect 13860 61852 13870 61908
rect 14130 61852 14140 61908
rect 14196 61852 14364 61908
rect 14420 61852 20412 61908
rect 20468 61852 20478 61908
rect 24882 61852 24892 61908
rect 24948 61852 25004 61908
rect 25060 61852 25070 61908
rect 2482 61740 2492 61796
rect 2548 61740 3164 61796
rect 3220 61740 3230 61796
rect 3714 61740 3724 61796
rect 3780 61740 5852 61796
rect 5908 61740 6972 61796
rect 7028 61740 7038 61796
rect 7196 61740 7756 61796
rect 7812 61740 7822 61796
rect 8418 61740 8428 61796
rect 8484 61740 10668 61796
rect 10724 61740 10734 61796
rect 12674 61740 12684 61796
rect 12740 61740 13356 61796
rect 13412 61740 13422 61796
rect 15698 61740 15708 61796
rect 15764 61740 21644 61796
rect 21700 61740 21710 61796
rect 22166 61740 22204 61796
rect 22260 61740 22270 61796
rect 26852 61740 29708 61796
rect 29764 61740 29774 61796
rect 3164 61684 3220 61740
rect 7196 61684 7252 61740
rect 2146 61628 2156 61684
rect 2212 61628 2380 61684
rect 2436 61628 2446 61684
rect 3164 61628 4172 61684
rect 4228 61628 4508 61684
rect 4564 61628 4574 61684
rect 6626 61628 6636 61684
rect 6692 61628 7196 61684
rect 7252 61628 7262 61684
rect 7522 61628 7532 61684
rect 7588 61628 9884 61684
rect 9940 61628 10780 61684
rect 10836 61628 10846 61684
rect 11340 61628 12628 61684
rect 13906 61628 13916 61684
rect 13972 61628 15036 61684
rect 15092 61628 15102 61684
rect 16930 61628 16940 61684
rect 16996 61628 21756 61684
rect 21812 61628 23772 61684
rect 23828 61628 23838 61684
rect 24182 61628 24220 61684
rect 24276 61628 24286 61684
rect 24546 61628 24556 61684
rect 24612 61628 25900 61684
rect 25956 61628 25966 61684
rect 2380 61460 2436 61628
rect 2706 61516 2716 61572
rect 2772 61516 4060 61572
rect 4116 61516 4126 61572
rect 5954 61516 5964 61572
rect 6020 61516 7420 61572
rect 7476 61516 7486 61572
rect 10210 61516 10220 61572
rect 10276 61516 10892 61572
rect 10948 61516 11116 61572
rect 11172 61516 11182 61572
rect 11340 61460 11396 61628
rect 12572 61572 12628 61628
rect 26852 61572 26908 61740
rect 12002 61516 12012 61572
rect 12068 61516 12348 61572
rect 12404 61516 12414 61572
rect 12572 61516 15148 61572
rect 15204 61516 15820 61572
rect 15876 61516 15886 61572
rect 18050 61516 18060 61572
rect 18116 61516 19740 61572
rect 19796 61516 26908 61572
rect 2380 61404 9100 61460
rect 9156 61404 9166 61460
rect 9874 61404 9884 61460
rect 9940 61404 11396 61460
rect 11890 61404 11900 61460
rect 11956 61404 14700 61460
rect 14756 61404 14924 61460
rect 14980 61404 14990 61460
rect 16034 61404 16044 61460
rect 16100 61404 16716 61460
rect 16772 61404 28028 61460
rect 28084 61404 29820 61460
rect 29876 61404 29886 61460
rect 1922 61292 1932 61348
rect 1988 61292 3612 61348
rect 3668 61292 6300 61348
rect 6356 61292 6366 61348
rect 7634 61292 7644 61348
rect 7700 61292 8428 61348
rect 8484 61292 8494 61348
rect 10658 61292 10668 61348
rect 10724 61292 12012 61348
rect 12068 61292 12078 61348
rect 13682 61292 13692 61348
rect 13748 61292 14028 61348
rect 14084 61292 14364 61348
rect 14420 61292 14430 61348
rect 14588 61292 15036 61348
rect 15092 61292 16940 61348
rect 16996 61292 17006 61348
rect 18162 61292 18172 61348
rect 18228 61292 20300 61348
rect 20356 61292 20366 61348
rect 21298 61292 21308 61348
rect 21364 61292 22652 61348
rect 22708 61292 22718 61348
rect 14588 61236 14644 61292
rect 20300 61236 20356 61292
rect 3154 61180 3164 61236
rect 3220 61180 4396 61236
rect 4452 61180 4956 61236
rect 5012 61180 5022 61236
rect 7298 61180 7308 61236
rect 7364 61180 8316 61236
rect 8372 61180 8382 61236
rect 13906 61180 13916 61236
rect 13972 61180 14644 61236
rect 14802 61180 14812 61236
rect 14868 61180 18844 61236
rect 18900 61180 18910 61236
rect 20300 61180 23100 61236
rect 23156 61180 23436 61236
rect 23492 61180 23502 61236
rect 30034 61180 30044 61236
rect 30100 61180 30110 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 5282 61068 5292 61124
rect 5348 61068 5852 61124
rect 5908 61068 6748 61124
rect 6804 61068 6814 61124
rect 8418 61068 8428 61124
rect 8484 61068 8652 61124
rect 8708 61068 8718 61124
rect 10098 61068 10108 61124
rect 10164 61068 14252 61124
rect 14308 61068 14318 61124
rect 14466 61068 14476 61124
rect 14532 61068 16828 61124
rect 16884 61068 16894 61124
rect 19142 61068 19180 61124
rect 19236 61068 19246 61124
rect 1922 60956 1932 61012
rect 1988 60956 3276 61012
rect 3332 60956 3342 61012
rect 4918 60956 4956 61012
rect 5012 60956 5022 61012
rect 6850 60956 6860 61012
rect 6916 60956 8988 61012
rect 9044 60956 9054 61012
rect 10182 60956 10220 61012
rect 10276 60956 10780 61012
rect 10836 60956 11116 61012
rect 11172 60956 11182 61012
rect 13682 60956 13692 61012
rect 13748 60956 16828 61012
rect 16884 60956 16894 61012
rect 18274 60956 18284 61012
rect 18340 60956 19068 61012
rect 19124 60956 19134 61012
rect 19730 60956 19740 61012
rect 19796 60956 22316 61012
rect 22372 60956 22382 61012
rect 3276 60900 3332 60956
rect 3276 60844 7644 60900
rect 7700 60844 7756 60900
rect 7812 60844 7822 60900
rect 13458 60844 13468 60900
rect 13524 60844 14028 60900
rect 14084 60844 14252 60900
rect 14308 60844 14318 60900
rect 14914 60844 14924 60900
rect 14980 60844 15820 60900
rect 15876 60844 16716 60900
rect 16772 60844 17612 60900
rect 17668 60844 17678 60900
rect 30044 60788 30100 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 3714 60732 3724 60788
rect 3780 60732 4172 60788
rect 4228 60732 4238 60788
rect 5478 60732 5516 60788
rect 5572 60732 5582 60788
rect 6262 60732 6300 60788
rect 6356 60732 6366 60788
rect 8642 60732 8652 60788
rect 8708 60732 9604 60788
rect 9762 60732 9772 60788
rect 9828 60732 14812 60788
rect 14868 60732 14878 60788
rect 15026 60732 15036 60788
rect 15092 60732 30100 60788
rect 9548 60676 9604 60732
rect 4050 60620 4060 60676
rect 4116 60620 7196 60676
rect 7252 60620 7262 60676
rect 8082 60620 8092 60676
rect 8148 60620 8652 60676
rect 8708 60620 8718 60676
rect 9548 60620 14476 60676
rect 14532 60620 14542 60676
rect 15698 60620 15708 60676
rect 15764 60620 16828 60676
rect 16884 60620 16894 60676
rect 20178 60620 20188 60676
rect 20244 60620 23212 60676
rect 23268 60620 23278 60676
rect 5170 60508 5180 60564
rect 5236 60508 7756 60564
rect 7812 60508 7822 60564
rect 8418 60508 8428 60564
rect 8484 60508 8988 60564
rect 9044 60508 9884 60564
rect 9940 60508 9950 60564
rect 10658 60508 10668 60564
rect 10724 60508 11900 60564
rect 11956 60508 11966 60564
rect 12338 60508 12348 60564
rect 12404 60508 12684 60564
rect 12740 60508 13020 60564
rect 13076 60508 13916 60564
rect 13972 60508 13982 60564
rect 16594 60508 16604 60564
rect 16660 60508 25340 60564
rect 25396 60508 25406 60564
rect 7858 60396 7868 60452
rect 7924 60396 11452 60452
rect 11508 60396 11518 60452
rect 11676 60396 12908 60452
rect 12964 60396 13692 60452
rect 13748 60396 13758 60452
rect 19142 60396 19180 60452
rect 19236 60396 19246 60452
rect 20850 60396 20860 60452
rect 20916 60396 22204 60452
rect 22260 60396 22270 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 11676 60340 11732 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 5730 60284 5740 60340
rect 5796 60284 11732 60340
rect 12114 60284 12124 60340
rect 12180 60284 16380 60340
rect 16436 60284 16446 60340
rect 26852 60284 30380 60340
rect 30436 60284 30446 60340
rect 26852 60228 26908 60284
rect 2594 60172 2604 60228
rect 2660 60172 6300 60228
rect 6356 60172 6366 60228
rect 7746 60172 7756 60228
rect 7812 60172 8204 60228
rect 8260 60172 8270 60228
rect 8530 60172 8540 60228
rect 8596 60172 8652 60228
rect 8708 60172 8718 60228
rect 9090 60172 9100 60228
rect 9156 60172 11228 60228
rect 11284 60172 11676 60228
rect 11732 60172 11742 60228
rect 12002 60172 12012 60228
rect 12068 60172 14140 60228
rect 14196 60172 14206 60228
rect 16258 60172 16268 60228
rect 16324 60172 20524 60228
rect 20580 60172 26908 60228
rect 27794 60172 27804 60228
rect 27860 60172 38108 60228
rect 38164 60172 38174 60228
rect 1586 60060 1596 60116
rect 1652 60060 3052 60116
rect 3108 60060 3118 60116
rect 4834 60060 4844 60116
rect 4900 60060 6188 60116
rect 6244 60060 6254 60116
rect 7522 60060 7532 60116
rect 7588 60060 8988 60116
rect 9044 60060 9054 60116
rect 9426 60060 9436 60116
rect 9492 60060 11564 60116
rect 11620 60060 11630 60116
rect 12786 60060 12796 60116
rect 12852 60060 13356 60116
rect 13412 60060 13422 60116
rect 14018 60060 14028 60116
rect 14084 60060 15820 60116
rect 15876 60060 15886 60116
rect 17826 60060 17836 60116
rect 17892 60060 18508 60116
rect 18564 60060 18574 60116
rect 23174 60060 23212 60116
rect 23268 60060 23278 60116
rect 15820 60004 15876 60060
rect 1250 59948 1260 60004
rect 1316 59948 4396 60004
rect 4452 59948 4462 60004
rect 6290 59948 6300 60004
rect 6356 59948 9772 60004
rect 9828 59948 9838 60004
rect 15820 59948 18284 60004
rect 18340 59948 18350 60004
rect 2482 59836 2492 59892
rect 2548 59836 4732 59892
rect 4788 59836 9996 59892
rect 10052 59836 10062 59892
rect 10220 59836 13580 59892
rect 13636 59836 13646 59892
rect 15362 59836 15372 59892
rect 15428 59836 19068 59892
rect 19124 59836 19134 59892
rect 4386 59724 4396 59780
rect 4452 59724 4844 59780
rect 4900 59724 4910 59780
rect 7074 59724 7084 59780
rect 7140 59724 8092 59780
rect 8148 59724 8158 59780
rect 10220 59668 10276 59836
rect 12674 59724 12684 59780
rect 12740 59724 12908 59780
rect 12964 59724 12974 59780
rect 17238 59724 17276 59780
rect 17332 59724 17342 59780
rect 17714 59724 17724 59780
rect 17780 59724 17948 59780
rect 18004 59724 18014 59780
rect 18172 59724 20860 59780
rect 20916 59724 20926 59780
rect 18172 59668 18228 59724
rect 5404 59612 10276 59668
rect 10546 59612 10556 59668
rect 10612 59612 12796 59668
rect 12852 59612 12862 59668
rect 13906 59612 13916 59668
rect 13972 59612 15932 59668
rect 15988 59612 18228 59668
rect 5404 59556 5460 59612
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 4732 59500 5460 59556
rect 5776 59500 5852 59556
rect 5908 59500 7644 59556
rect 7700 59500 7710 59556
rect 8642 59500 8652 59556
rect 8708 59500 11788 59556
rect 11844 59500 16604 59556
rect 16660 59500 16670 59556
rect 2818 59388 2828 59444
rect 2884 59388 3388 59444
rect 3444 59388 3454 59444
rect 4732 59332 4788 59500
rect 4946 59388 4956 59444
rect 5012 59388 7308 59444
rect 7364 59388 9100 59444
rect 9156 59388 9166 59444
rect 11218 59388 11228 59444
rect 11284 59388 11452 59444
rect 11508 59388 11518 59444
rect 15474 59388 15484 59444
rect 15540 59388 16268 59444
rect 16324 59388 16334 59444
rect 16930 59388 16940 59444
rect 16996 59388 21308 59444
rect 21364 59388 21374 59444
rect 3042 59276 3052 59332
rect 3108 59276 4788 59332
rect 8978 59276 8988 59332
rect 9044 59276 13580 59332
rect 13636 59276 13646 59332
rect 14130 59276 14140 59332
rect 14196 59276 18844 59332
rect 18900 59276 47852 59332
rect 47908 59276 47918 59332
rect 7942 59164 7980 59220
rect 8036 59164 8046 59220
rect 9762 59164 9772 59220
rect 9828 59164 9884 59220
rect 9940 59164 9950 59220
rect 10434 59164 10444 59220
rect 10500 59164 10556 59220
rect 10612 59164 10622 59220
rect 10994 59164 11004 59220
rect 11060 59164 18060 59220
rect 18116 59164 18126 59220
rect 4386 59052 4396 59108
rect 4452 59052 10220 59108
rect 10276 59052 10780 59108
rect 10836 59052 11340 59108
rect 11396 59052 11406 59108
rect 3266 58940 3276 58996
rect 3332 58940 3612 58996
rect 3668 58940 3678 58996
rect 4162 58940 4172 58996
rect 4228 58940 6076 58996
rect 6132 58940 6142 58996
rect 6290 58940 6300 58996
rect 6356 58940 10164 58996
rect 11442 58940 11452 58996
rect 11508 58940 15764 58996
rect 16818 58940 16828 58996
rect 16884 58940 16940 58996
rect 16996 58940 18172 58996
rect 18228 58940 19516 58996
rect 19572 58940 19582 58996
rect 10108 58884 10164 58940
rect 15708 58884 15764 58940
rect 6290 58828 6300 58884
rect 6356 58828 9604 58884
rect 10108 58828 14140 58884
rect 14196 58828 14206 58884
rect 15708 58828 19628 58884
rect 19684 58828 19694 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 9548 58772 9604 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 6290 58716 6300 58772
rect 6356 58716 6636 58772
rect 6692 58716 9324 58772
rect 9380 58716 9390 58772
rect 9548 58716 13804 58772
rect 13860 58716 13870 58772
rect 15026 58716 15036 58772
rect 15092 58716 15932 58772
rect 15988 58716 17724 58772
rect 17780 58716 17790 58772
rect 3714 58604 3724 58660
rect 3780 58604 15148 58660
rect 16594 58604 16604 58660
rect 16660 58604 16716 58660
rect 16772 58604 17164 58660
rect 17220 58604 17230 58660
rect 2594 58492 2604 58548
rect 2660 58492 5852 58548
rect 5908 58492 11564 58548
rect 11620 58492 11630 58548
rect 12114 58492 12124 58548
rect 12180 58492 12236 58548
rect 12292 58492 12302 58548
rect 12450 58492 12460 58548
rect 12516 58492 12572 58548
rect 12628 58492 12638 58548
rect 13654 58492 13692 58548
rect 13748 58492 13758 58548
rect 12460 58436 12516 58492
rect 3602 58380 3612 58436
rect 3668 58380 10332 58436
rect 10388 58380 10398 58436
rect 10658 58380 10668 58436
rect 10724 58380 12516 58436
rect 15092 58436 15148 58604
rect 15362 58492 15372 58548
rect 15428 58492 18956 58548
rect 19012 58492 19022 58548
rect 15092 58380 17500 58436
rect 17556 58380 17566 58436
rect 12460 58324 12516 58380
rect 5506 58268 5516 58324
rect 5572 58268 12292 58324
rect 12460 58268 22988 58324
rect 23044 58268 23054 58324
rect 12236 58212 12292 58268
rect 6402 58156 6412 58212
rect 6468 58156 6636 58212
rect 6692 58156 6702 58212
rect 7634 58156 7644 58212
rect 7700 58156 9548 58212
rect 9604 58156 12012 58212
rect 12068 58156 12078 58212
rect 12236 58156 14476 58212
rect 14532 58156 14542 58212
rect 19506 58156 19516 58212
rect 19572 58156 38668 58212
rect 38724 58156 38734 58212
rect 6178 58044 6188 58100
rect 6244 58044 6636 58100
rect 6692 58044 7196 58100
rect 7252 58044 7262 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 13804 57932 19180 57988
rect 19236 57932 19246 57988
rect 3378 57820 3388 57876
rect 3444 57820 7868 57876
rect 7924 57820 7934 57876
rect 8978 57820 8988 57876
rect 9044 57820 10780 57876
rect 10836 57820 10846 57876
rect 11554 57820 11564 57876
rect 11620 57820 12460 57876
rect 12516 57820 12526 57876
rect 13804 57764 13860 57932
rect 14690 57820 14700 57876
rect 14756 57820 15148 57876
rect 15204 57820 15214 57876
rect 2930 57708 2940 57764
rect 2996 57708 8764 57764
rect 8820 57708 13804 57764
rect 13860 57708 13870 57764
rect 12450 57596 12460 57652
rect 12516 57596 13804 57652
rect 13860 57596 13870 57652
rect 14242 57596 14252 57652
rect 14308 57596 15148 57652
rect 38658 57596 38668 57652
rect 38724 57596 40012 57652
rect 40068 57596 40078 57652
rect 15092 57540 15148 57596
rect 7298 57484 7308 57540
rect 7364 57484 10220 57540
rect 10276 57484 13356 57540
rect 13412 57484 14028 57540
rect 14084 57484 14700 57540
rect 14756 57484 14766 57540
rect 15092 57484 21308 57540
rect 21364 57484 21374 57540
rect 8082 57260 8092 57316
rect 8148 57260 13916 57316
rect 13972 57260 14252 57316
rect 14308 57260 14318 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 7858 57148 7868 57204
rect 7924 57148 10276 57204
rect 19478 57148 19516 57204
rect 19572 57148 19582 57204
rect 10220 57092 10276 57148
rect 8194 57036 8204 57092
rect 8260 57036 9996 57092
rect 10052 57036 10062 57092
rect 10220 57036 28476 57092
rect 28532 57036 28542 57092
rect 9202 56924 9212 56980
rect 9268 56924 9324 56980
rect 9380 56924 9390 56980
rect 9762 56924 9772 56980
rect 9828 56924 10108 56980
rect 10164 56924 10174 56980
rect 10332 56924 22540 56980
rect 22596 56924 22606 56980
rect 10332 56868 10388 56924
rect 4834 56812 4844 56868
rect 4900 56812 10388 56868
rect 13570 56812 13580 56868
rect 13636 56812 15148 56868
rect 15204 56812 15280 56868
rect 18396 56812 33180 56868
rect 33236 56812 33246 56868
rect 1586 56700 1596 56756
rect 1652 56700 3388 56756
rect 9314 56700 9324 56756
rect 9380 56700 18172 56756
rect 18228 56700 18238 56756
rect 3332 56196 3388 56700
rect 9762 56588 9772 56644
rect 9828 56588 11676 56644
rect 11732 56588 12908 56644
rect 12964 56588 12974 56644
rect 7970 56476 7980 56532
rect 8036 56476 12572 56532
rect 12628 56476 12638 56532
rect 12796 56476 17276 56532
rect 17332 56476 17342 56532
rect 12796 56308 12852 56476
rect 18396 56420 18452 56812
rect 18610 56588 18620 56644
rect 18676 56588 28812 56644
rect 28868 56588 28878 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 6402 56252 6412 56308
rect 6468 56252 12852 56308
rect 12908 56364 16380 56420
rect 16436 56364 18452 56420
rect 12908 56196 12964 56364
rect 14466 56252 14476 56308
rect 14532 56252 27804 56308
rect 27860 56252 27870 56308
rect 3332 56140 12964 56196
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 28802 55468 28812 55524
rect 28868 55468 29596 55524
rect 29652 55468 29662 55524
rect 21298 55356 21308 55412
rect 21364 55356 21868 55412
rect 21924 55356 21934 55412
rect 1362 55244 1372 55300
rect 1428 55244 8092 55300
rect 8148 55244 8158 55300
rect 10322 55244 10332 55300
rect 10388 55244 16828 55300
rect 16884 55244 16894 55300
rect 13906 55132 13916 55188
rect 13972 55132 25116 55188
rect 25172 55132 25182 55188
rect 4050 55020 4060 55076
rect 4116 55020 15708 55076
rect 15764 55020 15774 55076
rect 29922 55020 29932 55076
rect 29988 55020 77308 55076
rect 77364 55020 77374 55076
rect 3490 54908 3500 54964
rect 3556 54908 16156 54964
rect 16212 54908 16222 54964
rect 25106 54908 25116 54964
rect 25172 54908 26012 54964
rect 26068 54908 26078 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 3042 54796 3052 54852
rect 3108 54796 16492 54852
rect 16548 54796 16558 54852
rect 6626 54684 6636 54740
rect 6692 54684 40348 54740
rect 40404 54684 40414 54740
rect 2818 54460 2828 54516
rect 2884 54460 17724 54516
rect 17780 54460 17790 54516
rect 9650 54348 9660 54404
rect 9716 54348 27692 54404
rect 27748 54348 27758 54404
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 40338 53788 40348 53844
rect 40404 53788 41244 53844
rect 41300 53788 41310 53844
rect 7746 53676 7756 53732
rect 7812 53676 8316 53732
rect 8372 53676 25564 53732
rect 25620 53676 25630 53732
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 10322 51996 10332 52052
rect 10388 51996 36092 52052
rect 36148 51996 36158 52052
rect 6626 51884 6636 51940
rect 6692 51884 21420 51940
rect 21476 51884 21486 51940
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 11666 50316 11676 50372
rect 11732 50316 48860 50372
rect 48916 50316 48926 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 2706 49980 2716 50036
rect 2772 49980 21868 50036
rect 21924 49980 23212 50036
rect 23268 49980 23278 50036
rect 48850 49756 48860 49812
rect 48916 49756 49532 49812
rect 49588 49756 49598 49812
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 1474 48524 1484 48580
rect 1540 48524 19516 48580
rect 19572 48524 19582 48580
rect 9986 48300 9996 48356
rect 10052 48300 25676 48356
rect 25732 48300 25742 48356
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 7410 45164 7420 45220
rect 7476 45164 8204 45220
rect 8260 45164 13468 45220
rect 13524 45164 13534 45220
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 5954 43596 5964 43652
rect 6020 43596 17836 43652
rect 17892 43596 17902 43652
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 7522 41916 7532 41972
rect 7588 41916 32620 41972
rect 32676 41916 32686 41972
rect 4274 41804 4284 41860
rect 4340 41804 15148 41860
rect 15204 41804 15214 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 15138 40348 15148 40404
rect 15204 40348 15932 40404
rect 15988 40348 15998 40404
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 13794 36652 13804 36708
rect 13860 36652 17612 36708
rect 17668 36652 17678 36708
rect 17602 36204 17612 36260
rect 17668 36204 77420 36260
rect 77476 36204 77486 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 14802 6748 14812 6804
rect 14868 6748 17500 6804
rect 17556 6748 17566 6804
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 10994 6076 11004 6132
rect 11060 6076 12460 6132
rect 12516 6076 12526 6132
rect 49522 6076 49532 6132
rect 49588 6076 51212 6132
rect 51268 6076 52220 6132
rect 52276 6076 52286 6132
rect 8306 5964 8316 6020
rect 8372 5964 15036 6020
rect 15092 5964 15102 6020
rect 15922 5964 15932 6020
rect 15988 5964 18620 6020
rect 18676 5964 19628 6020
rect 19684 5964 19694 6020
rect 8194 5852 8204 5908
rect 8260 5852 52892 5908
rect 52948 5852 53340 5908
rect 53396 5852 53406 5908
rect 15362 5740 15372 5796
rect 15428 5740 18172 5796
rect 18228 5740 18844 5796
rect 18900 5740 18910 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 16706 5292 16716 5348
rect 16772 5292 46844 5348
rect 46900 5292 47740 5348
rect 47796 5292 47806 5348
rect 26002 5180 26012 5236
rect 26068 5180 34300 5236
rect 34356 5180 34748 5236
rect 34804 5180 34814 5236
rect 18834 5068 18844 5124
rect 18900 5068 22204 5124
rect 22260 5068 23436 5124
rect 23492 5068 26796 5124
rect 26852 5068 28028 5124
rect 28084 5068 32060 5124
rect 32116 5068 33292 5124
rect 33348 5068 34412 5124
rect 34468 5068 34972 5124
rect 35028 5068 39452 5124
rect 39508 5068 40684 5124
rect 40740 5068 47180 5124
rect 47236 5068 47964 5124
rect 48020 5068 51212 5124
rect 51268 5068 51772 5124
rect 51828 5068 51996 5124
rect 52052 5068 52332 5124
rect 52388 5068 53004 5124
rect 53060 5068 53070 5124
rect 24658 4844 24668 4900
rect 24724 4844 26012 4900
rect 26068 4844 26078 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 11218 4508 11228 4564
rect 11284 4508 11676 4564
rect 11732 4508 12348 4564
rect 12404 4508 14588 4564
rect 14644 4508 15372 4564
rect 15428 4508 15438 4564
rect 47842 4508 47852 4564
rect 47908 4508 50764 4564
rect 50820 4508 51772 4564
rect 51828 4508 51838 4564
rect 9986 4396 9996 4452
rect 10052 4396 11900 4452
rect 11956 4396 12796 4452
rect 12852 4396 12862 4452
rect 16594 4396 16604 4452
rect 16660 4396 17500 4452
rect 17556 4396 17566 4452
rect 19954 4396 19964 4452
rect 20020 4396 21420 4452
rect 21476 4396 21486 4452
rect 29586 4396 29596 4452
rect 29652 4396 30716 4452
rect 30772 4396 30782 4452
rect 35298 4396 35308 4452
rect 35364 4396 38332 4452
rect 38388 4396 38398 4452
rect 41010 4396 41020 4452
rect 41076 4396 43484 4452
rect 43540 4396 43550 4452
rect 48290 4396 48300 4452
rect 48356 4396 49532 4452
rect 49588 4396 49598 4452
rect 49858 4396 49868 4452
rect 49924 4396 50540 4452
rect 50596 4396 50606 4452
rect 52770 4396 52780 4452
rect 52836 4396 54908 4452
rect 54964 4396 54974 4452
rect 55234 4396 55244 4452
rect 55300 4396 55468 4452
rect 58258 4396 58268 4452
rect 58324 4396 64540 4452
rect 64596 4396 64606 4452
rect 66210 4396 66220 4452
rect 66276 4396 68460 4452
rect 68516 4396 68526 4452
rect 55412 4340 55468 4396
rect 7634 4284 7644 4340
rect 7700 4284 11340 4340
rect 11396 4284 11406 4340
rect 28354 4284 28364 4340
rect 28420 4284 29260 4340
rect 29316 4284 29326 4340
rect 53442 4284 53452 4340
rect 53508 4284 54012 4340
rect 54068 4284 54078 4340
rect 55412 4284 58604 4340
rect 58660 4284 58670 4340
rect 65314 4284 65324 4340
rect 65380 4284 65884 4340
rect 65940 4284 65950 4340
rect 74386 4284 74396 4340
rect 74452 4284 75180 4340
rect 75236 4284 77420 4340
rect 77476 4284 77486 4340
rect 52322 4172 52332 4228
rect 52388 4172 57932 4228
rect 57988 4172 57998 4228
rect 76066 4172 76076 4228
rect 76132 4172 77532 4228
rect 77588 4172 77598 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 6962 3612 6972 3668
rect 7028 3612 7868 3668
rect 7924 3612 7934 3668
rect 11666 3612 11676 3668
rect 11732 3612 12236 3668
rect 12292 3612 12302 3668
rect 15138 3612 15148 3668
rect 15204 3612 16044 3668
rect 16100 3612 16110 3668
rect 16370 3612 16380 3668
rect 16436 3612 18172 3668
rect 18228 3612 18238 3668
rect 21074 3612 21084 3668
rect 21140 3612 22092 3668
rect 22148 3612 22158 3668
rect 25778 3612 25788 3668
rect 25844 3612 26684 3668
rect 26740 3612 26750 3668
rect 30482 3612 30492 3668
rect 30548 3612 31388 3668
rect 31444 3612 31454 3668
rect 35186 3612 35196 3668
rect 35252 3612 35756 3668
rect 35812 3612 35822 3668
rect 39890 3612 39900 3668
rect 39956 3612 41692 3668
rect 41748 3612 41758 3668
rect 54002 3612 54012 3668
rect 54068 3612 54908 3668
rect 54964 3612 54974 3668
rect 58706 3612 58716 3668
rect 58772 3612 59276 3668
rect 59332 3612 59342 3668
rect 63410 3612 63420 3668
rect 63476 3612 65212 3668
rect 65268 3612 65278 3668
rect 68114 3612 68124 3668
rect 68180 3612 69132 3668
rect 69188 3612 69198 3668
rect 72818 3612 72828 3668
rect 72884 3612 73724 3668
rect 73780 3612 73790 3668
rect 1138 3500 1148 3556
rect 1204 3500 3500 3556
rect 3556 3500 4284 3556
rect 4340 3500 4350 3556
rect 38658 3500 38668 3556
rect 38724 3500 41020 3556
rect 41076 3500 41086 3556
rect 41234 3500 41244 3556
rect 41300 3500 51660 3556
rect 51716 3500 52780 3556
rect 52836 3500 52846 3556
rect 53330 3500 53340 3556
rect 53396 3500 65324 3556
rect 65380 3500 65390 3556
rect 72594 3500 72604 3556
rect 72660 3500 73276 3556
rect 73332 3500 77308 3556
rect 77364 3500 77374 3556
rect 44604 3388 45612 3444
rect 45668 3388 45678 3444
rect 44604 3332 44660 3388
rect 44594 3276 44604 3332
rect 44660 3276 44670 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 21532 79212 21588 79268
rect 17612 78204 17668 78260
rect 6748 78092 6804 78148
rect 4956 77980 5012 78036
rect 4284 77756 4340 77812
rect 7308 77644 7364 77700
rect 7644 77532 7700 77588
rect 24220 77308 24276 77364
rect 3500 77196 3556 77252
rect 3276 76860 3332 76916
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 33292 76748 33348 76804
rect 6524 76524 6580 76580
rect 21420 76300 21476 76356
rect 11004 76188 11060 76244
rect 30604 76188 30660 76244
rect 3836 75964 3892 76020
rect 9996 76076 10052 76132
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 9884 75964 9940 76020
rect 2044 75852 2100 75908
rect 6972 75852 7028 75908
rect 9212 75740 9268 75796
rect 14140 75740 14196 75796
rect 4172 75628 4228 75684
rect 26124 75628 26180 75684
rect 7532 75516 7588 75572
rect 17724 75516 17780 75572
rect 4060 75404 4116 75460
rect 4844 75404 4900 75460
rect 13468 75404 13524 75460
rect 22988 75404 23044 75460
rect 3052 75180 3108 75236
rect 3500 75180 3556 75236
rect 10780 75292 10836 75348
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 5740 75068 5796 75124
rect 29596 75068 29652 75124
rect 33628 75068 33684 75124
rect 15148 74956 15204 75012
rect 30604 74956 30660 75012
rect 9772 74844 9828 74900
rect 12684 74844 12740 74900
rect 2604 74732 2660 74788
rect 11788 74732 11844 74788
rect 25564 74732 25620 74788
rect 7420 74620 7476 74676
rect 10332 74620 10388 74676
rect 1260 74508 1316 74564
rect 5516 74508 5572 74564
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 32060 74508 32116 74564
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 3388 74284 3444 74340
rect 4060 74284 4116 74340
rect 13468 74284 13524 74340
rect 12684 74172 12740 74228
rect 31612 74172 31668 74228
rect 2156 74060 2212 74116
rect 15148 74060 15204 74116
rect 3500 73948 3556 74004
rect 3948 73948 4004 74004
rect 6860 73948 6916 74004
rect 7756 73948 7812 74004
rect 8092 73948 8148 74004
rect 9660 73948 9716 74004
rect 10444 73948 10500 74004
rect 16156 73948 16212 74004
rect 21644 73948 21700 74004
rect 29596 73948 29652 74004
rect 31612 73948 31668 74004
rect 33628 73948 33684 74004
rect 5964 73836 6020 73892
rect 6412 73836 6468 73892
rect 7196 73836 7252 73892
rect 32956 73836 33012 73892
rect 4172 73724 4228 73780
rect 5292 73724 5348 73780
rect 8092 73724 8148 73780
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 1372 73612 1428 73668
rect 8540 73612 8596 73668
rect 6076 73388 6132 73444
rect 10668 73388 10724 73444
rect 2044 73276 2100 73332
rect 5180 73276 5236 73332
rect 6188 73276 6244 73332
rect 8316 73276 8372 73332
rect 17724 73276 17780 73332
rect 2940 73164 2996 73220
rect 4060 73164 4116 73220
rect 7756 73164 7812 73220
rect 10444 73164 10500 73220
rect 20188 73164 20244 73220
rect 25340 73164 25396 73220
rect 27804 73164 27860 73220
rect 5068 73052 5124 73108
rect 29820 73052 29876 73108
rect 8540 72940 8596 72996
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 6636 72828 6692 72884
rect 6076 72716 6132 72772
rect 10668 72716 10724 72772
rect 10892 72716 10948 72772
rect 19516 72716 19572 72772
rect 2044 72604 2100 72660
rect 7196 72604 7252 72660
rect 29820 72604 29876 72660
rect 1484 72492 1540 72548
rect 5068 72492 5124 72548
rect 7084 72492 7140 72548
rect 12236 72492 12292 72548
rect 8540 72380 8596 72436
rect 10220 72380 10276 72436
rect 16380 72380 16436 72436
rect 23996 72380 24052 72436
rect 24444 72380 24500 72436
rect 5628 72268 5684 72324
rect 5852 72268 5908 72324
rect 9996 72268 10052 72324
rect 19516 72268 19572 72324
rect 32172 72268 32228 72324
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 7532 72044 7588 72100
rect 10108 72044 10164 72100
rect 12796 72044 12852 72100
rect 16156 71932 16212 71988
rect 5740 71820 5796 71876
rect 5964 71820 6020 71876
rect 10220 71820 10276 71876
rect 2380 71708 2436 71764
rect 3276 71708 3332 71764
rect 4172 71708 4228 71764
rect 5516 71708 5572 71764
rect 1596 71596 1652 71652
rect 8540 71596 8596 71652
rect 32956 71484 33012 71540
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 8092 71260 8148 71316
rect 29596 71148 29652 71204
rect 4284 71036 4340 71092
rect 8652 71036 8708 71092
rect 3276 70924 3332 70980
rect 4956 70924 5012 70980
rect 6300 70924 6356 70980
rect 6524 70924 6580 70980
rect 25452 70812 25508 70868
rect 23996 70700 24052 70756
rect 32172 70700 32228 70756
rect 33292 70700 33348 70756
rect 5180 70588 5236 70644
rect 6860 70588 6916 70644
rect 10556 70588 10612 70644
rect 12348 70588 12404 70644
rect 21308 70588 21364 70644
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 5964 70476 6020 70532
rect 27356 70476 27412 70532
rect 32172 70476 32228 70532
rect 32620 70476 32676 70532
rect 2716 70364 2772 70420
rect 5740 70364 5796 70420
rect 6076 70364 6132 70420
rect 6748 70364 6804 70420
rect 7532 70364 7588 70420
rect 8092 70364 8148 70420
rect 10444 70252 10500 70308
rect 11452 70252 11508 70308
rect 18732 70252 18788 70308
rect 3724 70140 3780 70196
rect 11788 70140 11844 70196
rect 16604 70140 16660 70196
rect 17836 70140 17892 70196
rect 32508 70140 32564 70196
rect 7308 70028 7364 70084
rect 8652 70028 8708 70084
rect 9436 70028 9492 70084
rect 13468 70028 13524 70084
rect 25676 70028 25732 70084
rect 27356 70028 27412 70084
rect 5628 69916 5684 69972
rect 11116 69804 11172 69860
rect 11452 69804 11508 69860
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 9324 69692 9380 69748
rect 3836 69580 3892 69636
rect 7196 69580 7252 69636
rect 7980 69580 8036 69636
rect 18508 69580 18564 69636
rect 28588 69580 28644 69636
rect 9548 69468 9604 69524
rect 32508 69468 32564 69524
rect 7644 69356 7700 69412
rect 9324 69356 9380 69412
rect 11900 69356 11956 69412
rect 5740 69244 5796 69300
rect 6076 69244 6132 69300
rect 9996 69244 10052 69300
rect 11676 69244 11732 69300
rect 7196 69132 7252 69188
rect 9884 69132 9940 69188
rect 18060 69020 18116 69076
rect 28588 69132 28644 69188
rect 31724 69132 31780 69188
rect 21756 69020 21812 69076
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4284 68908 4340 68964
rect 4956 68908 5012 68964
rect 3164 68796 3220 68852
rect 15484 68796 15540 68852
rect 2828 68684 2884 68740
rect 3948 68684 4004 68740
rect 17500 68684 17556 68740
rect 21868 68572 21924 68628
rect 6972 68460 7028 68516
rect 8428 68460 8484 68516
rect 10444 68460 10500 68516
rect 21756 68460 21812 68516
rect 1148 68348 1204 68404
rect 5292 68348 5348 68404
rect 11004 68348 11060 68404
rect 22316 68572 22372 68628
rect 24892 68572 24948 68628
rect 4956 68236 5012 68292
rect 16940 68236 16996 68292
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 3836 68124 3892 68180
rect 15148 68124 15204 68180
rect 9436 68012 9492 68068
rect 10444 68012 10500 68068
rect 18284 68012 18340 68068
rect 9324 67900 9380 67956
rect 4284 67788 4340 67844
rect 15036 67788 15092 67844
rect 22092 67788 22148 67844
rect 24220 67788 24276 67844
rect 17500 67676 17556 67732
rect 22316 67676 22372 67732
rect 3276 67564 3332 67620
rect 5068 67564 5124 67620
rect 21980 67564 22036 67620
rect 27580 67564 27636 67620
rect 24444 67452 24500 67508
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 2380 67340 2436 67396
rect 3276 67340 3332 67396
rect 9324 67340 9380 67396
rect 15596 67340 15652 67396
rect 6748 67228 6804 67284
rect 7868 67228 7924 67284
rect 10444 67228 10500 67284
rect 12796 67228 12852 67284
rect 15036 67228 15092 67284
rect 18060 67116 18116 67172
rect 26124 67116 26180 67172
rect 4956 67004 5012 67060
rect 15260 67004 15316 67060
rect 15484 67004 15540 67060
rect 16604 67004 16660 67060
rect 4284 66892 4340 66948
rect 6748 66892 6804 66948
rect 10668 66892 10724 66948
rect 12012 66892 12068 66948
rect 14252 66892 14308 66948
rect 16940 66892 16996 66948
rect 17948 66892 18004 66948
rect 7644 66780 7700 66836
rect 7868 66780 7924 66836
rect 8764 66780 8820 66836
rect 18284 66780 18340 66836
rect 27580 66780 27636 66836
rect 4956 66668 5012 66724
rect 9436 66668 9492 66724
rect 9884 66668 9940 66724
rect 14028 66668 14084 66724
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 5180 66556 5236 66612
rect 5964 66556 6020 66612
rect 7756 66556 7812 66612
rect 11116 66556 11172 66612
rect 24780 66556 24836 66612
rect 6636 66444 6692 66500
rect 26124 66444 26180 66500
rect 13692 66332 13748 66388
rect 6636 66220 6692 66276
rect 7196 66220 7252 66276
rect 9100 66220 9156 66276
rect 9436 66108 9492 66164
rect 11676 66108 11732 66164
rect 22316 66108 22372 66164
rect 6636 65996 6692 66052
rect 14028 65996 14084 66052
rect 22204 65996 22260 66052
rect 3612 65884 3668 65940
rect 4956 65884 5012 65940
rect 8316 65884 8372 65940
rect 8764 65884 8820 65940
rect 11676 65884 11732 65940
rect 15260 65884 15316 65940
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 3724 65772 3780 65828
rect 7196 65660 7252 65716
rect 7980 65660 8036 65716
rect 8316 65660 8372 65716
rect 12460 65660 12516 65716
rect 17500 65660 17556 65716
rect 18172 65660 18228 65716
rect 25452 65660 25508 65716
rect 26684 65660 26740 65716
rect 22540 65548 22596 65604
rect 11452 65436 11508 65492
rect 16828 65436 16884 65492
rect 3052 65324 3108 65380
rect 13916 65324 13972 65380
rect 15596 65324 15652 65380
rect 16492 65324 16548 65380
rect 20188 65324 20244 65380
rect 3836 65212 3892 65268
rect 4844 65212 4900 65268
rect 10108 65212 10164 65268
rect 16268 65212 16324 65268
rect 18508 65212 18564 65268
rect 3724 65100 3780 65156
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 6636 64988 6692 65044
rect 18396 64988 18452 65044
rect 12460 64876 12516 64932
rect 12908 64876 12964 64932
rect 14028 64876 14084 64932
rect 8540 64764 8596 64820
rect 10220 64764 10276 64820
rect 15484 64764 15540 64820
rect 15820 64764 15876 64820
rect 3276 64652 3332 64708
rect 7196 64652 7252 64708
rect 18732 64652 18788 64708
rect 3052 64540 3108 64596
rect 4956 64540 5012 64596
rect 7868 64428 7924 64484
rect 12236 64428 12292 64484
rect 6972 64316 7028 64372
rect 10444 64316 10500 64372
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 15484 64204 15540 64260
rect 19628 64204 19684 64260
rect 26684 64204 26740 64260
rect 4956 64092 5012 64148
rect 12236 64092 12292 64148
rect 14028 64092 14084 64148
rect 3836 63980 3892 64036
rect 8652 63980 8708 64036
rect 3276 63868 3332 63924
rect 18396 63868 18452 63924
rect 18732 63868 18788 63924
rect 19628 63868 19684 63924
rect 26684 63868 26740 63924
rect 7084 63756 7140 63812
rect 10220 63756 10276 63812
rect 17612 63756 17668 63812
rect 26908 63756 26964 63812
rect 2380 63644 2436 63700
rect 7308 63532 7364 63588
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 2716 63420 2772 63476
rect 3612 63308 3668 63364
rect 7980 63308 8036 63364
rect 11564 63308 11620 63364
rect 16716 63308 16772 63364
rect 14028 63196 14084 63252
rect 6188 63084 6244 63140
rect 4284 62972 4340 63028
rect 13580 62972 13636 63028
rect 7756 62860 7812 62916
rect 4844 62636 4900 62692
rect 11900 62636 11956 62692
rect 23212 62860 23268 62916
rect 22092 62748 22148 62804
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 21532 62524 21588 62580
rect 3164 62412 3220 62468
rect 12236 62412 12292 62468
rect 17276 62412 17332 62468
rect 21980 62412 22036 62468
rect 5292 62300 5348 62356
rect 3388 62188 3444 62244
rect 3948 62188 4004 62244
rect 24780 62188 24836 62244
rect 5068 62076 5124 62132
rect 9996 62076 10052 62132
rect 12012 62076 12068 62132
rect 15708 62076 15764 62132
rect 18732 61964 18788 62020
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 7532 61852 7588 61908
rect 24892 61852 24948 61908
rect 10668 61740 10724 61796
rect 21644 61740 21700 61796
rect 22204 61740 22260 61796
rect 2156 61628 2212 61684
rect 24220 61628 24276 61684
rect 7420 61516 7476 61572
rect 10892 61516 10948 61572
rect 9100 61404 9156 61460
rect 10668 61292 10724 61348
rect 14028 61292 14084 61348
rect 15036 61292 15092 61348
rect 14812 61180 14868 61236
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 8428 61068 8484 61124
rect 14476 61068 14532 61124
rect 16828 61068 16884 61124
rect 19180 61068 19236 61124
rect 4956 60956 5012 61012
rect 10220 60956 10276 61012
rect 7644 60844 7700 60900
rect 16716 60844 16772 60900
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4172 60732 4228 60788
rect 5516 60732 5572 60788
rect 6300 60732 6356 60788
rect 14812 60732 14868 60788
rect 8652 60620 8708 60676
rect 14476 60620 14532 60676
rect 15708 60620 15764 60676
rect 5180 60508 5236 60564
rect 16604 60508 16660 60564
rect 25340 60508 25396 60564
rect 12908 60396 12964 60452
rect 13692 60396 13748 60452
rect 19180 60396 19236 60452
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 5740 60284 5796 60340
rect 6300 60172 6356 60228
rect 8540 60172 8596 60228
rect 27804 60172 27860 60228
rect 4844 60060 4900 60116
rect 7532 60060 7588 60116
rect 14028 60060 14084 60116
rect 23212 60060 23268 60116
rect 1260 59948 1316 60004
rect 9772 59948 9828 60004
rect 13580 59836 13636 59892
rect 12684 59724 12740 59780
rect 17276 59724 17332 59780
rect 17948 59724 18004 59780
rect 13916 59612 13972 59668
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 5852 59500 5908 59556
rect 11788 59500 11844 59556
rect 16604 59500 16660 59556
rect 2828 59388 2884 59444
rect 16268 59388 16324 59444
rect 14140 59276 14196 59332
rect 7980 59164 8036 59220
rect 9884 59164 9940 59220
rect 10556 59164 10612 59220
rect 11004 59164 11060 59220
rect 3276 58940 3332 58996
rect 3612 58940 3668 58996
rect 16940 58940 16996 58996
rect 6300 58828 6356 58884
rect 14140 58828 14196 58884
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 13804 58716 13860 58772
rect 15036 58716 15092 58772
rect 16604 58604 16660 58660
rect 2604 58492 2660 58548
rect 11564 58492 11620 58548
rect 12236 58492 12292 58548
rect 12460 58492 12516 58548
rect 13692 58492 13748 58548
rect 3612 58380 3668 58436
rect 10332 58380 10388 58436
rect 5516 58268 5572 58324
rect 22988 58268 23044 58324
rect 6412 58156 6468 58212
rect 9548 58156 9604 58212
rect 19516 58156 19572 58212
rect 6188 58044 6244 58100
rect 6636 58044 6692 58100
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 10780 57820 10836 57876
rect 13804 57596 13860 57652
rect 21308 57484 21364 57540
rect 13916 57260 13972 57316
rect 14252 57260 14308 57316
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 7868 57148 7924 57204
rect 19516 57148 19572 57204
rect 9212 56924 9268 56980
rect 10108 56924 10164 56980
rect 22540 56924 22596 56980
rect 15148 56812 15204 56868
rect 1596 56700 1652 56756
rect 18172 56700 18228 56756
rect 9772 56588 9828 56644
rect 17276 56476 17332 56532
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 16380 56364 16436 56420
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 21308 55356 21364 55412
rect 1372 55244 1428 55300
rect 10332 55244 10388 55300
rect 13916 55132 13972 55188
rect 4060 55020 4116 55076
rect 3500 54908 3556 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 3052 54796 3108 54852
rect 16492 54796 16548 54852
rect 6636 54684 6692 54740
rect 17724 54460 17780 54516
rect 9660 54348 9716 54404
rect 27692 54348 27748 54404
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 25564 53676 25620 53732
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 21420 51884 21476 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 1484 48524 1540 48580
rect 25676 48300 25732 48356
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 13468 45164 13524 45220
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 17836 43596 17892 43652
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 7532 41916 7588 41972
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 1148 3500 1204 3556
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 21532 79268 21588 79278
rect 17612 78260 17668 78270
rect 6748 78148 6804 78158
rect 4956 78036 5012 78046
rect 4284 77812 4340 77822
rect 3500 77252 3556 77262
rect 3276 76916 3332 76926
rect 2044 75908 2100 75918
rect 1260 74564 1316 74574
rect 1148 68404 1204 68414
rect 1148 3556 1204 68348
rect 1260 60004 1316 74508
rect 1260 59938 1316 59948
rect 1372 73668 1428 73678
rect 1372 55300 1428 73612
rect 2044 73332 2100 75852
rect 3052 75236 3108 75246
rect 2604 74788 2660 74798
rect 2044 72660 2100 73276
rect 2044 72594 2100 72604
rect 2156 74116 2212 74126
rect 1372 55234 1428 55244
rect 1484 72548 1540 72558
rect 1484 48580 1540 72492
rect 1596 71652 1652 71662
rect 1596 56756 1652 71596
rect 2156 61684 2212 74060
rect 2380 71764 2436 71774
rect 2380 67396 2436 71708
rect 2380 63700 2436 67340
rect 2380 63634 2436 63644
rect 2156 61618 2212 61628
rect 2604 58548 2660 74732
rect 2940 73220 2996 73230
rect 2716 70420 2772 70430
rect 2716 63476 2772 70364
rect 2716 63410 2772 63420
rect 2828 68740 2884 68750
rect 2828 59444 2884 68684
rect 2828 59378 2884 59388
rect 2604 58482 2660 58492
rect 1596 56690 1652 56700
rect 2940 55468 2996 73164
rect 3052 65380 3108 75180
rect 3276 71764 3332 76860
rect 3500 75236 3556 77196
rect 3500 75170 3556 75180
rect 3836 76020 3892 76030
rect 3276 71698 3332 71708
rect 3388 74340 3444 74350
rect 3276 70980 3332 70990
rect 3052 64596 3108 65324
rect 3052 64530 3108 64540
rect 3164 68852 3220 68862
rect 3164 62468 3220 68796
rect 3276 67620 3332 70924
rect 3276 67554 3332 67564
rect 3276 67396 3332 67406
rect 3276 64708 3332 67340
rect 3276 64642 3332 64652
rect 3164 62402 3220 62412
rect 3276 63924 3332 63934
rect 3276 58996 3332 63868
rect 3388 62244 3444 74284
rect 3388 62178 3444 62188
rect 3500 74004 3556 74014
rect 3276 58930 3332 58940
rect 2940 55412 3108 55468
rect 3052 54852 3108 55412
rect 3500 54964 3556 73948
rect 3724 70196 3780 70206
rect 3612 65940 3668 65950
rect 3612 63364 3668 65884
rect 3724 65828 3780 70140
rect 3836 69636 3892 75964
rect 4172 75684 4228 75694
rect 4060 75460 4116 75470
rect 4060 74340 4116 75404
rect 4060 74274 4116 74284
rect 3836 69570 3892 69580
rect 3948 74004 4004 74014
rect 3948 68964 4004 73948
rect 4172 73780 4228 75628
rect 4172 73714 4228 73724
rect 3836 68908 4004 68964
rect 4060 73220 4116 73230
rect 3836 68180 3892 68908
rect 3836 68114 3892 68124
rect 3948 68740 4004 68750
rect 3724 65156 3780 65772
rect 3724 65090 3780 65100
rect 3836 65268 3892 65278
rect 3836 64036 3892 65212
rect 3836 63970 3892 63980
rect 3612 63298 3668 63308
rect 3948 62244 4004 68684
rect 3948 62178 4004 62188
rect 3612 58996 3668 59006
rect 3612 58436 3668 58940
rect 3612 58370 3668 58380
rect 4060 55076 4116 73164
rect 4172 71764 4228 71774
rect 4172 60788 4228 71708
rect 4284 71092 4340 77756
rect 4284 71026 4340 71036
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4284 68964 4340 68974
rect 4284 67844 4340 68908
rect 4284 67778 4340 67788
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4284 66948 4340 66958
rect 4284 63028 4340 66892
rect 4284 62962 4340 62972
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4844 75460 4900 75470
rect 4844 65268 4900 75404
rect 4956 70980 5012 77980
rect 6524 76580 6580 76590
rect 5740 75124 5796 75134
rect 5516 74564 5572 74574
rect 5292 73780 5348 73790
rect 5180 73332 5236 73342
rect 5068 73108 5124 73118
rect 5068 72548 5124 73052
rect 5068 72482 5124 72492
rect 4956 70914 5012 70924
rect 5180 70644 5236 73276
rect 5180 70578 5236 70588
rect 4956 68964 5012 68974
rect 4956 68292 5012 68908
rect 4956 68226 5012 68236
rect 5292 68404 5348 73724
rect 5068 67620 5124 67630
rect 4956 67060 5012 67070
rect 4956 66724 5012 67004
rect 4956 66658 5012 66668
rect 4844 65202 4900 65212
rect 4956 65940 5012 65950
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4956 64596 5012 65884
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4172 60722 4228 60732
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4060 55010 4116 55020
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4844 64540 4956 64596
rect 4844 62692 4900 64540
rect 4956 64530 5012 64540
rect 4844 60116 4900 62636
rect 4956 64148 5012 64158
rect 4956 61012 5012 64092
rect 5068 62132 5124 67564
rect 5068 62066 5124 62076
rect 5180 66612 5236 66622
rect 4956 60946 5012 60956
rect 5180 60564 5236 66556
rect 5292 62356 5348 68348
rect 5292 62290 5348 62300
rect 5516 71764 5572 74508
rect 5180 60498 5236 60508
rect 5516 60788 5572 71708
rect 5628 72324 5684 72334
rect 5628 69972 5684 72268
rect 5740 71876 5796 75068
rect 5964 73892 6020 73902
rect 5740 70420 5796 71820
rect 5740 70354 5796 70364
rect 5852 72324 5908 72334
rect 5628 69906 5684 69916
rect 4844 60050 4900 60060
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 5516 58324 5572 60732
rect 5740 69300 5796 69310
rect 5740 60340 5796 69244
rect 5740 60274 5796 60284
rect 5852 59556 5908 72268
rect 5964 71876 6020 73836
rect 6412 73892 6468 73902
rect 6076 73444 6132 73454
rect 6076 72772 6132 73388
rect 6076 72706 6132 72716
rect 6188 73332 6244 73342
rect 5964 71810 6020 71820
rect 5964 70532 6020 70542
rect 5964 66612 6020 70476
rect 6076 70420 6132 70430
rect 6076 69300 6132 70364
rect 6076 69234 6132 69244
rect 5964 66546 6020 66556
rect 5852 59490 5908 59500
rect 6188 63140 6244 73276
rect 5516 58258 5572 58268
rect 6188 58100 6244 63084
rect 6300 70980 6356 70990
rect 6300 60788 6356 70924
rect 6300 60228 6356 60732
rect 6300 58884 6356 60172
rect 6300 58818 6356 58828
rect 6412 58212 6468 73836
rect 6524 70980 6580 76524
rect 6524 70914 6580 70924
rect 6636 72884 6692 72894
rect 6636 66500 6692 72828
rect 6748 70420 6804 78092
rect 7308 77700 7364 77710
rect 6972 75908 7028 75918
rect 6860 74004 6916 74014
rect 6860 70644 6916 73948
rect 6860 70578 6916 70588
rect 6748 70354 6804 70364
rect 6972 68516 7028 75852
rect 7196 73892 7252 73902
rect 7196 72660 7252 73836
rect 6748 67284 6804 67294
rect 6748 66948 6804 67228
rect 6748 66882 6804 66892
rect 6636 66276 6692 66444
rect 6636 66210 6692 66220
rect 6636 66052 6692 66062
rect 6636 65044 6692 65996
rect 6636 64978 6692 64988
rect 6972 64372 7028 68460
rect 6972 64306 7028 64316
rect 7084 72548 7140 72558
rect 7084 63812 7140 72492
rect 7196 69636 7252 72604
rect 7308 70084 7364 77644
rect 7644 77588 7700 77598
rect 7532 75572 7588 75582
rect 7308 70018 7364 70028
rect 7420 74676 7476 74686
rect 7196 69570 7252 69580
rect 7196 69188 7252 69198
rect 7196 66276 7252 69132
rect 7252 66220 7364 66276
rect 7196 66210 7252 66220
rect 7084 63746 7140 63756
rect 7196 65716 7252 65726
rect 7196 64708 7252 65660
rect 6412 58146 6468 58156
rect 6188 58034 6244 58044
rect 6636 58100 6692 58110
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 3500 54898 3556 54908
rect 3052 54786 3108 54796
rect 1484 48514 1540 48524
rect 4448 54124 4768 55636
rect 6636 54740 6692 58044
rect 6636 54674 6692 54684
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 7196 50428 7252 64652
rect 7308 63588 7364 66220
rect 7308 63522 7364 63532
rect 7420 61572 7476 74620
rect 7532 72100 7588 75516
rect 7532 72034 7588 72044
rect 7420 61506 7476 61516
rect 7532 70420 7588 70430
rect 7532 61908 7588 70364
rect 7532 60116 7588 61852
rect 7644 69412 7700 77532
rect 11004 76244 11060 76254
rect 9996 76132 10052 76142
rect 9884 76020 9940 76030
rect 9212 75796 9268 75806
rect 7756 74004 7812 74014
rect 7756 73220 7812 73948
rect 8092 74004 8148 74014
rect 8092 73780 8148 73948
rect 8092 73714 8148 73724
rect 8540 73668 8596 73678
rect 7756 73154 7812 73164
rect 8316 73332 8372 73342
rect 8092 71316 8148 71326
rect 8092 70420 8148 71260
rect 8092 70354 8148 70364
rect 7644 66836 7700 69356
rect 7980 69636 8036 69646
rect 7644 60900 7700 66780
rect 7868 67284 7924 67294
rect 7868 66836 7924 67228
rect 7868 66770 7924 66780
rect 7756 66612 7812 66622
rect 7756 62916 7812 66556
rect 7980 65716 8036 69580
rect 7980 65650 8036 65660
rect 8316 65940 8372 73276
rect 8540 72996 8596 73612
rect 8540 72930 8596 72940
rect 8540 72436 8596 72446
rect 8540 71652 8596 72380
rect 8540 71586 8596 71596
rect 8652 71092 8708 71102
rect 8652 70084 8708 71036
rect 8316 65716 8372 65884
rect 8316 65650 8372 65660
rect 8428 68516 8484 68526
rect 7756 62850 7812 62860
rect 7868 64484 7924 64494
rect 7644 60834 7700 60844
rect 7532 60050 7588 60060
rect 7868 57204 7924 64428
rect 7980 63364 8036 63374
rect 7980 59220 8036 63308
rect 8428 61124 8484 68460
rect 8428 61058 8484 61068
rect 8540 64820 8596 64830
rect 8540 60228 8596 64764
rect 8652 64036 8708 70028
rect 8764 66836 8820 66846
rect 8764 65940 8820 66780
rect 8764 65874 8820 65884
rect 9100 66276 9156 66286
rect 8652 60676 8708 63980
rect 9100 61460 9156 66220
rect 9100 61394 9156 61404
rect 8652 60610 8708 60620
rect 8540 60162 8596 60172
rect 7980 59154 8036 59164
rect 7868 57138 7924 57148
rect 9212 56980 9268 75740
rect 9772 74900 9828 74910
rect 9660 74004 9716 74014
rect 9436 70084 9492 70094
rect 9324 69748 9380 69758
rect 9324 69412 9380 69692
rect 9324 69346 9380 69356
rect 9436 68068 9492 70028
rect 9436 68002 9492 68012
rect 9548 69524 9604 69534
rect 9324 67956 9380 67966
rect 9324 67396 9380 67900
rect 9324 67330 9380 67340
rect 9436 66724 9492 66734
rect 9436 66164 9492 66668
rect 9436 66098 9492 66108
rect 9548 58212 9604 69468
rect 9548 58146 9604 58156
rect 9212 56914 9268 56924
rect 9660 54404 9716 73948
rect 9772 60004 9828 74844
rect 9884 69188 9940 75964
rect 9996 72324 10052 76076
rect 10780 75348 10836 75358
rect 10332 74676 10388 74686
rect 9996 72258 10052 72268
rect 10220 72436 10276 72446
rect 10108 72100 10164 72110
rect 9884 69122 9940 69132
rect 9996 69300 10052 69310
rect 9772 56644 9828 59948
rect 9884 66724 9940 66734
rect 9884 59220 9940 66668
rect 9996 62132 10052 69244
rect 9996 62066 10052 62076
rect 10108 65268 10164 72044
rect 9884 59154 9940 59164
rect 10108 56980 10164 65212
rect 10220 71876 10276 72380
rect 10220 64820 10276 71820
rect 10220 64754 10276 64764
rect 10220 63812 10276 63822
rect 10220 61012 10276 63756
rect 10220 60946 10276 60956
rect 10108 56914 10164 56924
rect 10332 58436 10388 74620
rect 10444 74004 10500 74014
rect 10444 73220 10500 73948
rect 10444 70308 10500 73164
rect 10668 73444 10724 73454
rect 10668 72772 10724 73388
rect 10668 72706 10724 72716
rect 10444 70242 10500 70252
rect 10556 70644 10612 70654
rect 10444 68516 10500 68526
rect 10444 68068 10500 68460
rect 10444 68002 10500 68012
rect 10444 67284 10500 67294
rect 10444 64372 10500 67228
rect 10444 64306 10500 64316
rect 10556 59220 10612 70588
rect 10668 66948 10724 66958
rect 10668 61796 10724 66892
rect 10668 61348 10724 61740
rect 10668 61282 10724 61292
rect 10556 59154 10612 59164
rect 9772 56578 9828 56588
rect 10332 55300 10388 58380
rect 10780 57876 10836 75292
rect 10892 72772 10948 72782
rect 10892 61572 10948 72716
rect 10892 61506 10948 61516
rect 11004 68404 11060 76188
rect 14140 75796 14196 75806
rect 13468 75460 13524 75470
rect 12684 74900 12740 74910
rect 11788 74788 11844 74798
rect 11452 70308 11508 70318
rect 11004 59220 11060 68348
rect 11116 69860 11172 69870
rect 11116 66612 11172 69804
rect 11116 66546 11172 66556
rect 11452 69860 11508 70252
rect 11452 65492 11508 69804
rect 11788 70196 11844 74732
rect 12684 74228 12740 74844
rect 11676 69300 11732 69310
rect 11676 66164 11732 69244
rect 11676 65940 11732 66108
rect 11676 65874 11732 65884
rect 11452 65426 11508 65436
rect 11004 59154 11060 59164
rect 11564 63364 11620 63374
rect 11564 58548 11620 63308
rect 11788 59556 11844 70140
rect 12236 72548 12292 72558
rect 11900 69412 11956 69422
rect 11900 62692 11956 69356
rect 11900 62626 11956 62636
rect 12012 66948 12068 66958
rect 12012 62132 12068 66892
rect 12236 64484 12292 72492
rect 12236 64148 12292 64428
rect 12236 64082 12292 64092
rect 12348 70644 12404 70654
rect 12012 62066 12068 62076
rect 12236 62468 12292 62478
rect 12348 62468 12404 70588
rect 12292 62412 12404 62468
rect 12460 65716 12516 65726
rect 12460 64932 12516 65660
rect 11788 59490 11844 59500
rect 11564 58482 11620 58492
rect 12236 58548 12292 62412
rect 12236 58482 12292 58492
rect 12460 58548 12516 64876
rect 12684 59780 12740 74172
rect 13468 74340 13524 75404
rect 12796 72100 12852 72110
rect 12796 67284 12852 72044
rect 12796 67218 12852 67228
rect 13468 70084 13524 74284
rect 12908 64932 12964 64942
rect 12908 60452 12964 64876
rect 12908 60386 12964 60396
rect 12684 59714 12740 59724
rect 12460 58482 12516 58492
rect 10780 57810 10836 57820
rect 10332 55234 10388 55244
rect 9660 54338 9716 54348
rect 7196 50372 7588 50428
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 1148 3490 1204 3500
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 7532 41972 7588 50372
rect 13468 45220 13524 70028
rect 14028 66724 14084 66734
rect 13692 66388 13748 66398
rect 13580 63028 13636 63038
rect 13580 59892 13636 62972
rect 13692 62188 13748 66332
rect 14028 66052 14084 66668
rect 13916 65380 13972 65390
rect 13692 62132 13860 62188
rect 13580 59826 13636 59836
rect 13692 60452 13748 60462
rect 13692 58548 13748 60396
rect 13692 58482 13748 58492
rect 13804 58772 13860 62132
rect 13916 59668 13972 65324
rect 14028 64932 14084 65996
rect 14028 64866 14084 64876
rect 14028 64148 14084 64158
rect 14028 63252 14084 64092
rect 14028 61348 14084 63196
rect 14028 60116 14084 61292
rect 14028 60050 14084 60060
rect 13916 59602 13972 59612
rect 14140 59332 14196 75740
rect 15148 75012 15204 75022
rect 15148 74116 15204 74956
rect 15148 68180 15204 74060
rect 16156 74004 16212 74014
rect 16156 71988 16212 73948
rect 16156 71922 16212 71932
rect 16380 72436 16436 72446
rect 15036 67844 15092 67854
rect 15036 67284 15092 67788
rect 15036 67218 15092 67228
rect 14140 58884 14196 59276
rect 14140 58818 14196 58828
rect 14252 66948 14308 66958
rect 13804 57652 13860 58716
rect 13804 57586 13860 57596
rect 13916 57316 13972 57326
rect 13916 55188 13972 57260
rect 14252 57316 14308 66892
rect 15036 61348 15092 61358
rect 14812 61236 14868 61246
rect 14476 61124 14532 61134
rect 14476 60676 14532 61068
rect 14812 60788 14868 61180
rect 14812 60722 14868 60732
rect 14476 60610 14532 60620
rect 15036 58772 15092 61292
rect 15036 58706 15092 58716
rect 14252 57250 14308 57260
rect 15148 56868 15204 68124
rect 15484 68852 15540 68862
rect 15260 67060 15316 67070
rect 15260 65940 15316 67004
rect 15484 67060 15540 68796
rect 15484 66994 15540 67004
rect 15596 67396 15652 67406
rect 15260 65874 15316 65884
rect 15596 65380 15652 67340
rect 15596 65314 15652 65324
rect 16268 65268 16324 65278
rect 15484 64820 15540 64830
rect 15484 64260 15540 64764
rect 15484 64194 15540 64204
rect 15820 64820 15876 64830
rect 15820 63028 15876 64764
rect 15708 62972 15876 63028
rect 15708 62132 15764 62972
rect 15708 60676 15764 62076
rect 15708 60610 15764 60620
rect 16268 59444 16324 65212
rect 16268 59378 16324 59388
rect 15148 56802 15204 56812
rect 16380 56420 16436 72380
rect 16604 70196 16660 70206
rect 16604 67060 16660 70140
rect 17500 68740 17556 68750
rect 16604 66994 16660 67004
rect 16940 68292 16996 68302
rect 16940 66948 16996 68236
rect 16828 65492 16884 65502
rect 16380 56354 16436 56364
rect 16492 65380 16548 65390
rect 13916 55122 13972 55132
rect 16492 54852 16548 65324
rect 16716 63364 16772 63374
rect 16716 60900 16772 63308
rect 16828 61124 16884 65436
rect 16828 61058 16884 61068
rect 16716 60834 16772 60844
rect 16604 60564 16660 60574
rect 16604 59556 16660 60508
rect 16604 58660 16660 59500
rect 16940 58996 16996 66892
rect 17500 67732 17556 68684
rect 17500 65716 17556 67676
rect 17500 65650 17556 65660
rect 17612 63812 17668 78204
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 17612 63746 17668 63756
rect 17724 75572 17780 75582
rect 17724 73332 17780 75516
rect 16940 58930 16996 58940
rect 17276 62468 17332 62478
rect 17276 59780 17332 62412
rect 16604 58594 16660 58604
rect 17276 56532 17332 59724
rect 17276 56466 17332 56476
rect 16492 54786 16548 54796
rect 17724 54516 17780 73276
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19516 72772 19572 72782
rect 19516 72324 19572 72716
rect 18732 70308 18788 70318
rect 17724 54450 17780 54460
rect 17836 70196 17892 70206
rect 13468 45154 13524 45164
rect 17836 43652 17892 70140
rect 18508 69636 18564 69646
rect 18060 69076 18116 69086
rect 18060 67172 18116 69020
rect 18060 67106 18116 67116
rect 18284 68068 18340 68078
rect 17948 66948 18004 66958
rect 17948 59780 18004 66892
rect 18284 66836 18340 68012
rect 18284 66770 18340 66780
rect 17948 59714 18004 59724
rect 18172 65716 18228 65726
rect 18172 56756 18228 65660
rect 18508 65268 18564 69580
rect 18508 65202 18564 65212
rect 18396 65044 18452 65054
rect 18396 63924 18452 64988
rect 18732 64708 18788 70252
rect 18732 64642 18788 64652
rect 18396 63858 18452 63868
rect 18732 63924 18788 63934
rect 18732 62020 18788 63868
rect 18732 61954 18788 61964
rect 19180 61124 19236 61134
rect 19180 60452 19236 61068
rect 19180 60386 19236 60396
rect 19516 58212 19572 72268
rect 19808 72156 20128 73668
rect 21420 76356 21476 76366
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 20188 73220 20244 73230
rect 20188 65380 20244 73164
rect 20188 65314 20244 65324
rect 21308 70644 21364 70654
rect 19628 64260 19684 64270
rect 19628 63924 19684 64204
rect 19628 63858 19684 63868
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19516 57204 19572 58156
rect 19516 57138 19572 57148
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 18172 56690 18228 56700
rect 17836 43586 17892 43596
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 21308 57540 21364 70588
rect 21308 55412 21364 57484
rect 21308 55346 21364 55356
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 21420 51940 21476 76300
rect 21532 62580 21588 79212
rect 24220 77364 24276 77374
rect 22988 75460 23044 75470
rect 21532 62514 21588 62524
rect 21644 74004 21700 74014
rect 21644 61796 21700 73948
rect 21756 69076 21812 69086
rect 21756 68516 21812 69020
rect 21868 68628 21924 68638
rect 22316 68628 22372 68638
rect 21924 68572 22316 68628
rect 21868 68562 21924 68572
rect 22316 68562 22372 68572
rect 21756 68450 21812 68460
rect 22092 67844 22148 67854
rect 21980 67620 22036 67630
rect 21980 62468 22036 67564
rect 22092 62804 22148 67788
rect 22316 67732 22372 67742
rect 22316 66164 22372 67676
rect 22316 66098 22372 66108
rect 22092 62738 22148 62748
rect 22204 66052 22260 66062
rect 21980 62402 22036 62412
rect 21644 61730 21700 61740
rect 22204 61796 22260 65996
rect 22204 61730 22260 61740
rect 22540 65604 22596 65614
rect 22540 56980 22596 65548
rect 22988 58324 23044 75404
rect 23996 72436 24052 72446
rect 23996 70756 24052 72380
rect 23996 70690 24052 70700
rect 24220 67844 24276 77308
rect 33292 76804 33348 76814
rect 30604 76244 30660 76254
rect 26124 75684 26180 75694
rect 25564 74788 25620 74798
rect 25340 73220 25396 73230
rect 23212 62916 23268 62926
rect 23212 60116 23268 62860
rect 24220 61684 24276 67788
rect 24444 72436 24500 72446
rect 24444 67508 24500 72380
rect 24444 67442 24500 67452
rect 24892 68628 24948 68638
rect 24780 66612 24836 66622
rect 24780 62244 24836 66556
rect 24780 62178 24836 62188
rect 24892 61908 24948 68572
rect 24892 61842 24948 61852
rect 24220 61618 24276 61628
rect 25340 60564 25396 73164
rect 25452 70868 25508 70878
rect 25452 65716 25508 70812
rect 25452 65650 25508 65660
rect 25340 60498 25396 60508
rect 23212 60050 23268 60060
rect 22988 58258 23044 58268
rect 22540 56914 22596 56924
rect 25564 53732 25620 74732
rect 25564 53666 25620 53676
rect 25676 70084 25732 70094
rect 21420 51874 21476 51884
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 25676 48356 25732 70028
rect 26124 67172 26180 75628
rect 29596 75124 29652 75134
rect 29596 74004 29652 75068
rect 30604 75012 30660 76188
rect 30604 74946 30660 74956
rect 32060 74564 32116 74574
rect 27804 73220 27860 73230
rect 27356 70532 27412 70542
rect 27356 70084 27412 70476
rect 27356 70018 27412 70028
rect 26124 66500 26180 67116
rect 27580 67620 27636 67630
rect 27580 66836 27636 67564
rect 27580 66770 27636 66780
rect 26124 66434 26180 66444
rect 26684 65716 26740 65726
rect 26684 65604 26740 65660
rect 26684 65548 26964 65604
rect 26684 64260 26740 64270
rect 26684 63924 26740 64204
rect 26684 63858 26740 63868
rect 26908 63812 26964 65548
rect 26908 63746 26964 63756
rect 27804 60228 27860 73164
rect 29596 71204 29652 73948
rect 31612 74228 31668 74238
rect 31612 74004 31668 74172
rect 31612 73938 31668 73948
rect 29820 73108 29876 73118
rect 29820 72660 29876 73052
rect 29820 72594 29876 72604
rect 29596 71138 29652 71148
rect 32060 70588 32116 74508
rect 32956 73892 33012 73902
rect 32172 72324 32228 72334
rect 32172 70756 32228 72268
rect 32956 71540 33012 73836
rect 32956 71474 33012 71484
rect 32172 70690 32228 70700
rect 33292 70756 33348 76748
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 33628 75124 33684 75134
rect 33628 74004 33684 75068
rect 33628 73938 33684 73948
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 33292 70690 33348 70700
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 31724 70532 32116 70588
rect 32172 70532 32228 70542
rect 32620 70532 32676 70542
rect 28588 69636 28644 69646
rect 28588 69188 28644 69580
rect 28588 69122 28644 69132
rect 31724 69188 31780 70532
rect 32228 70476 32620 70532
rect 32172 70466 32228 70476
rect 32620 70466 32676 70476
rect 32508 70196 32564 70206
rect 32508 69524 32564 70140
rect 32508 69458 32564 69468
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 31724 69122 31780 69132
rect 27804 55468 27860 60172
rect 27692 55412 27860 55468
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 27692 54404 27748 55412
rect 27692 54338 27748 54348
rect 25676 48290 25732 48300
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 7532 41906 7588 41916
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__I gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6944 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A1
timestamp 1669390400
transform 1 0 7280 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A2
timestamp 1669390400
transform 1 0 6720 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__I
timestamp 1669390400
transform 1 0 16912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__A1
timestamp 1669390400
transform -1 0 5376 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__A2
timestamp 1669390400
transform -1 0 2464 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1669390400
transform -1 0 4256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I
timestamp 1669390400
transform -1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A1
timestamp 1669390400
transform 1 0 12768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A2
timestamp 1669390400
transform 1 0 12320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A1
timestamp 1669390400
transform 1 0 12432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A2
timestamp 1669390400
transform -1 0 12208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__A1
timestamp 1669390400
transform -1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__A2
timestamp 1669390400
transform 1 0 14560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A1
timestamp 1669390400
transform 1 0 19600 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A2
timestamp 1669390400
transform -1 0 18256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A1
timestamp 1669390400
transform -1 0 22848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A2
timestamp 1669390400
transform 1 0 22176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A1
timestamp 1669390400
transform 1 0 27216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A2
timestamp 1669390400
transform 1 0 26768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A1
timestamp 1669390400
transform -1 0 32704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A2
timestamp 1669390400
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__A1
timestamp 1669390400
transform -1 0 34384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__A2
timestamp 1669390400
transform -1 0 34384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A1
timestamp 1669390400
transform -1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A2
timestamp 1669390400
transform 1 0 39424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__A1
timestamp 1669390400
transform -1 0 46928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__A2
timestamp 1669390400
transform 1 0 47152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__A1
timestamp 1669390400
transform 1 0 53312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__A2
timestamp 1669390400
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__A1
timestamp 1669390400
transform 1 0 51184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__A2
timestamp 1669390400
transform -1 0 51856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A1
timestamp 1669390400
transform 1 0 50736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A2
timestamp 1669390400
transform 1 0 51184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A1
timestamp 1669390400
transform -1 0 51744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A2
timestamp 1669390400
transform -1 0 52192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__I
timestamp 1669390400
transform 1 0 65296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A1
timestamp 1669390400
transform 1 0 17584 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A2
timestamp 1669390400
transform 1 0 18032 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__I
timestamp 1669390400
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__I
timestamp 1669390400
transform -1 0 10752 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__A1
timestamp 1669390400
transform 1 0 27552 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__A2
timestamp 1669390400
transform 1 0 28784 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1669390400
transform 1 0 30912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A2
timestamp 1669390400
transform -1 0 29904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__I
timestamp 1669390400
transform -1 0 2800 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__I
timestamp 1669390400
transform -1 0 11312 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A1
timestamp 1669390400
transform -1 0 4704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A2
timestamp 1669390400
transform -1 0 2016 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__288__I
timestamp 1669390400
transform -1 0 2240 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__I
timestamp 1669390400
transform 1 0 21504 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A1
timestamp 1669390400
transform 1 0 21728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1669390400
transform -1 0 24304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__B1
timestamp 1669390400
transform 1 0 22624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__B2
timestamp 1669390400
transform -1 0 22400 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__A1
timestamp 1669390400
transform -1 0 3584 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A1
timestamp 1669390400
transform 1 0 35504 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A2
timestamp 1669390400
transform 1 0 31360 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A3
timestamp 1669390400
transform -1 0 35280 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__A4
timestamp 1669390400
transform 1 0 34608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A1
timestamp 1669390400
transform -1 0 2016 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A2
timestamp 1669390400
transform -1 0 2688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A3
timestamp 1669390400
transform -1 0 3024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A4
timestamp 1669390400
transform -1 0 2464 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A1
timestamp 1669390400
transform -1 0 35728 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A2
timestamp 1669390400
transform 1 0 35056 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A3
timestamp 1669390400
transform 1 0 35504 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A4
timestamp 1669390400
transform 1 0 35952 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A1
timestamp 1669390400
transform 1 0 36288 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A2
timestamp 1669390400
transform 1 0 34944 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A3
timestamp 1669390400
transform 1 0 35840 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A4
timestamp 1669390400
transform 1 0 35392 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A1
timestamp 1669390400
transform 1 0 39872 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A4
timestamp 1669390400
transform 1 0 39424 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A1
timestamp 1669390400
transform 1 0 6272 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A2
timestamp 1669390400
transform -1 0 4592 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A1
timestamp 1669390400
transform -1 0 17808 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A2
timestamp 1669390400
transform -1 0 20720 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A3
timestamp 1669390400
transform -1 0 20272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A4
timestamp 1669390400
transform -1 0 19600 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A1
timestamp 1669390400
transform 1 0 11872 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A2
timestamp 1669390400
transform 1 0 11424 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__I
timestamp 1669390400
transform -1 0 6832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A1
timestamp 1669390400
transform -1 0 2688 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A2
timestamp 1669390400
transform -1 0 2464 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A3
timestamp 1669390400
transform 1 0 2912 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A4
timestamp 1669390400
transform -1 0 2128 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A1
timestamp 1669390400
transform -1 0 4704 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A2
timestamp 1669390400
transform -1 0 4256 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A3
timestamp 1669390400
transform -1 0 4256 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A1
timestamp 1669390400
transform 1 0 4928 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A2
timestamp 1669390400
transform 1 0 5824 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A3
timestamp 1669390400
transform 1 0 5712 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A4
timestamp 1669390400
transform -1 0 6384 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A1
timestamp 1669390400
transform 1 0 15120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1669390400
transform 1 0 16688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A1
timestamp 1669390400
transform -1 0 4032 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A2
timestamp 1669390400
transform -1 0 5936 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A3
timestamp 1669390400
transform -1 0 3136 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A4
timestamp 1669390400
transform -1 0 3808 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__A1
timestamp 1669390400
transform 1 0 21056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__A2
timestamp 1669390400
transform -1 0 23408 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__B1
timestamp 1669390400
transform 1 0 22736 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__307__B2
timestamp 1669390400
transform 1 0 20384 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__I
timestamp 1669390400
transform -1 0 6160 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__I
timestamp 1669390400
transform -1 0 12656 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A1
timestamp 1669390400
transform -1 0 13664 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A2
timestamp 1669390400
transform 1 0 10752 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__B
timestamp 1669390400
transform -1 0 12208 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A1
timestamp 1669390400
transform 1 0 8064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A2
timestamp 1669390400
transform 1 0 8960 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A3
timestamp 1669390400
transform 1 0 3136 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A1
timestamp 1669390400
transform -1 0 11200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A2
timestamp 1669390400
transform -1 0 10304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__A1
timestamp 1669390400
transform 1 0 6720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__A2
timestamp 1669390400
transform 1 0 4928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__B1
timestamp 1669390400
transform 1 0 4032 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__B2
timestamp 1669390400
transform -1 0 3808 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__A1
timestamp 1669390400
transform 1 0 7168 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A1
timestamp 1669390400
transform -1 0 2688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A2
timestamp 1669390400
transform -1 0 4032 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A1
timestamp 1669390400
transform 1 0 6272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A2
timestamp 1669390400
transform 1 0 7056 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A3
timestamp 1669390400
transform 1 0 5824 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A4
timestamp 1669390400
transform 1 0 3584 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__317__A1
timestamp 1669390400
transform 1 0 3136 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__A1
timestamp 1669390400
transform -1 0 5936 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__A1
timestamp 1669390400
transform 1 0 7616 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A1
timestamp 1669390400
transform 1 0 6608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A3
timestamp 1669390400
transform -1 0 7392 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__A1
timestamp 1669390400
transform 1 0 4480 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__A2
timestamp 1669390400
transform 1 0 4928 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A1
timestamp 1669390400
transform -1 0 2016 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A2
timestamp 1669390400
transform -1 0 2240 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__B
timestamp 1669390400
transform -1 0 3024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__A1
timestamp 1669390400
transform 1 0 2688 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__A1
timestamp 1669390400
transform 1 0 2688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__A2
timestamp 1669390400
transform 1 0 3136 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__B
timestamp 1669390400
transform -1 0 2016 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__A1
timestamp 1669390400
transform 1 0 2688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__A2
timestamp 1669390400
transform 1 0 4480 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__I
timestamp 1669390400
transform -1 0 13776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A1
timestamp 1669390400
transform 1 0 4032 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__A2
timestamp 1669390400
transform -1 0 4256 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__B
timestamp 1669390400
transform -1 0 5600 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A1
timestamp 1669390400
transform 1 0 14448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A2
timestamp 1669390400
transform 1 0 14224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A3
timestamp 1669390400
transform 1 0 13552 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__A4
timestamp 1669390400
transform -1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__A1
timestamp 1669390400
transform -1 0 4144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__A3
timestamp 1669390400
transform -1 0 2016 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__A1
timestamp 1669390400
transform 1 0 3584 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__A2
timestamp 1669390400
transform 1 0 4032 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A1
timestamp 1669390400
transform -1 0 1904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__A2
timestamp 1669390400
transform -1 0 7840 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__A1
timestamp 1669390400
transform 1 0 4928 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A1
timestamp 1669390400
transform 1 0 38752 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A2
timestamp 1669390400
transform 1 0 38304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__A3
timestamp 1669390400
transform 1 0 39872 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__A1
timestamp 1669390400
transform 1 0 8064 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__B
timestamp 1669390400
transform 1 0 8064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A1
timestamp 1669390400
transform 1 0 10192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__A2
timestamp 1669390400
transform -1 0 9968 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__A1
timestamp 1669390400
transform -1 0 3920 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__A2
timestamp 1669390400
transform -1 0 4368 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__A1
timestamp 1669390400
transform 1 0 36400 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__A2
timestamp 1669390400
transform 1 0 29792 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__A1
timestamp 1669390400
transform 1 0 18480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__A3
timestamp 1669390400
transform 1 0 19824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__A1
timestamp 1669390400
transform 1 0 17136 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__A2
timestamp 1669390400
transform -1 0 18256 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__A1
timestamp 1669390400
transform -1 0 8736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__A2
timestamp 1669390400
transform -1 0 2464 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__A1
timestamp 1669390400
transform -1 0 9408 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__A2
timestamp 1669390400
transform -1 0 9856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__A3
timestamp 1669390400
transform 1 0 2688 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A1
timestamp 1669390400
transform 1 0 6720 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A2
timestamp 1669390400
transform 1 0 9968 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__B
timestamp 1669390400
transform 1 0 3136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A1
timestamp 1669390400
transform -1 0 2016 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__A2
timestamp 1669390400
transform 1 0 4704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__B
timestamp 1669390400
transform -1 0 2464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__I
timestamp 1669390400
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__A1
timestamp 1669390400
transform 1 0 3584 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__A2
timestamp 1669390400
transform -1 0 9856 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__B
timestamp 1669390400
transform -1 0 6384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A1
timestamp 1669390400
transform 1 0 12880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A2
timestamp 1669390400
transform 1 0 6272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A3
timestamp 1669390400
transform -1 0 2016 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A1
timestamp 1669390400
transform 1 0 4928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A3
timestamp 1669390400
transform 1 0 5824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__A1
timestamp 1669390400
transform 1 0 18704 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__A2
timestamp 1669390400
transform 1 0 18256 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__B
timestamp 1669390400
transform 1 0 19152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__A1
timestamp 1669390400
transform 1 0 4480 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__A2
timestamp 1669390400
transform -1 0 3696 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__B
timestamp 1669390400
transform -1 0 4144 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A1
timestamp 1669390400
transform 1 0 6272 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__A2
timestamp 1669390400
transform -1 0 6944 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__B
timestamp 1669390400
transform 1 0 7168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A1
timestamp 1669390400
transform -1 0 2464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A2
timestamp 1669390400
transform -1 0 3360 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__A3
timestamp 1669390400
transform 1 0 3584 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A1
timestamp 1669390400
transform 1 0 3584 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A2
timestamp 1669390400
transform -1 0 3472 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A3
timestamp 1669390400
transform -1 0 2464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__A1
timestamp 1669390400
transform -1 0 3808 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__A2
timestamp 1669390400
transform -1 0 4928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A1
timestamp 1669390400
transform 1 0 6832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A2
timestamp 1669390400
transform -1 0 7840 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__A1
timestamp 1669390400
transform 1 0 10752 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__A2
timestamp 1669390400
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A1
timestamp 1669390400
transform 1 0 16240 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A2
timestamp 1669390400
transform 1 0 14336 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__A1
timestamp 1669390400
transform -1 0 19824 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__A2
timestamp 1669390400
transform 1 0 17584 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__B1
timestamp 1669390400
transform -1 0 16912 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__B2
timestamp 1669390400
transform 1 0 10864 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1669390400
transform 1 0 20048 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1669390400
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A2
timestamp 1669390400
transform 1 0 27664 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1669390400
transform -1 0 2576 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A2
timestamp 1669390400
transform -1 0 3472 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__B1
timestamp 1669390400
transform -1 0 3584 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__B2
timestamp 1669390400
transform -1 0 2128 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A1
timestamp 1669390400
transform -1 0 2912 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A2
timestamp 1669390400
transform -1 0 3808 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A1
timestamp 1669390400
transform 1 0 5824 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A2
timestamp 1669390400
transform 1 0 4928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A3
timestamp 1669390400
transform 1 0 8400 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A1
timestamp 1669390400
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A2
timestamp 1669390400
transform -1 0 28560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1669390400
transform -1 0 2016 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A2
timestamp 1669390400
transform -1 0 9072 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__B1
timestamp 1669390400
transform 1 0 7616 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__B2
timestamp 1669390400
transform -1 0 8400 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__C
timestamp 1669390400
transform 1 0 8736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A1
timestamp 1669390400
transform 1 0 18704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__A2
timestamp 1669390400
transform 1 0 19152 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__B1
timestamp 1669390400
transform -1 0 19824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__B2
timestamp 1669390400
transform -1 0 17136 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A1
timestamp 1669390400
transform -1 0 4256 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A2
timestamp 1669390400
transform 1 0 4928 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I
timestamp 1669390400
transform -1 0 6496 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A1
timestamp 1669390400
transform 1 0 7168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A2
timestamp 1669390400
transform -1 0 6048 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__A1
timestamp 1669390400
transform -1 0 4704 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__A2
timestamp 1669390400
transform -1 0 5600 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1669390400
transform 1 0 10640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A2
timestamp 1669390400
transform 1 0 11200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__I0
timestamp 1669390400
transform 1 0 8848 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__374__S
timestamp 1669390400
transform 1 0 12992 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__A1
timestamp 1669390400
transform -1 0 4480 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__A2
timestamp 1669390400
transform -1 0 2912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__B1
timestamp 1669390400
transform 1 0 3360 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__B2
timestamp 1669390400
transform -1 0 5936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__C
timestamp 1669390400
transform -1 0 2464 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A1
timestamp 1669390400
transform -1 0 16016 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__377__A2
timestamp 1669390400
transform -1 0 14224 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A1
timestamp 1669390400
transform 1 0 8176 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A2
timestamp 1669390400
transform 1 0 8624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A1
timestamp 1669390400
transform 1 0 7168 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A2
timestamp 1669390400
transform 1 0 7728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__A1
timestamp 1669390400
transform 1 0 9296 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__381__A2
timestamp 1669390400
transform -1 0 7952 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__A1
timestamp 1669390400
transform 1 0 3360 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__383__A2
timestamp 1669390400
transform -1 0 3136 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1669390400
transform -1 0 10528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A2
timestamp 1669390400
transform 1 0 13776 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__B1
timestamp 1669390400
transform -1 0 12656 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__B2
timestamp 1669390400
transform -1 0 13104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__C1
timestamp 1669390400
transform -1 0 12096 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__C2
timestamp 1669390400
transform -1 0 2464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__A1
timestamp 1669390400
transform -1 0 5600 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__385__A2
timestamp 1669390400
transform -1 0 6608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A1
timestamp 1669390400
transform -1 0 14784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2
timestamp 1669390400
transform 1 0 13552 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1669390400
transform 1 0 7168 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A2
timestamp 1669390400
transform 1 0 7616 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__A1
timestamp 1669390400
transform -1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A1
timestamp 1669390400
transform 1 0 3024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A2
timestamp 1669390400
transform -1 0 2688 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1669390400
transform 1 0 12320 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A2
timestamp 1669390400
transform 1 0 14448 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__B
timestamp 1669390400
transform 1 0 11984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A1
timestamp 1669390400
transform -1 0 14336 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1669390400
transform 1 0 11536 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__B1
timestamp 1669390400
transform 1 0 9968 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__B2
timestamp 1669390400
transform -1 0 15120 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A1
timestamp 1669390400
transform 1 0 15232 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A2
timestamp 1669390400
transform 1 0 17136 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A1
timestamp 1669390400
transform 1 0 12656 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A2
timestamp 1669390400
transform 1 0 14672 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1669390400
transform 1 0 14000 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A2
timestamp 1669390400
transform 1 0 12768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1
timestamp 1669390400
transform 1 0 11424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1669390400
transform 1 0 15344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A1
timestamp 1669390400
transform 1 0 33488 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A2
timestamp 1669390400
transform 1 0 33936 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A1
timestamp 1669390400
transform 1 0 37744 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__A2
timestamp 1669390400
transform 1 0 35952 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__B1
timestamp 1669390400
transform 1 0 36400 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__B2
timestamp 1669390400
transform -1 0 19936 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__C
timestamp 1669390400
transform 1 0 38192 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A1
timestamp 1669390400
transform 1 0 34608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__A2
timestamp 1669390400
transform 1 0 34160 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A1
timestamp 1669390400
transform -1 0 15456 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A2
timestamp 1669390400
transform -1 0 15904 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__A1
timestamp 1669390400
transform 1 0 19712 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__A2
timestamp 1669390400
transform 1 0 19264 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1669390400
transform 1 0 15792 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1669390400
transform -1 0 17360 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__B
timestamp 1669390400
transform 1 0 12880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A1
timestamp 1669390400
transform -1 0 2912 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__A2
timestamp 1669390400
transform -1 0 3920 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__B
timestamp 1669390400
transform -1 0 3360 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A1
timestamp 1669390400
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__A2
timestamp 1669390400
transform 1 0 26320 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__B
timestamp 1669390400
transform 1 0 26768 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A1
timestamp 1669390400
transform 1 0 19488 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A2
timestamp 1669390400
transform 1 0 34832 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__B1
timestamp 1669390400
transform 1 0 22736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__B2
timestamp 1669390400
transform -1 0 21840 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A1
timestamp 1669390400
transform 1 0 35280 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A1
timestamp 1669390400
transform -1 0 12544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A2
timestamp 1669390400
transform -1 0 11312 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A2
timestamp 1669390400
transform -1 0 9072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A4
timestamp 1669390400
transform -1 0 15008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A1
timestamp 1669390400
transform -1 0 16464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__A2
timestamp 1669390400
transform -1 0 16576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__C
timestamp 1669390400
transform 1 0 17584 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A1
timestamp 1669390400
transform -1 0 19152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A2
timestamp 1669390400
transform -1 0 18368 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1669390400
transform 1 0 20832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A2
timestamp 1669390400
transform 1 0 20608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1669390400
transform 1 0 36848 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A2
timestamp 1669390400
transform 1 0 37408 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__B1
timestamp 1669390400
transform 1 0 37744 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__B2
timestamp 1669390400
transform 1 0 36400 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__C1
timestamp 1669390400
transform -1 0 21840 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__C2
timestamp 1669390400
transform 1 0 37296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A1
timestamp 1669390400
transform 1 0 39088 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1669390400
transform -1 0 17808 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1669390400
transform 1 0 41440 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__B
timestamp 1669390400
transform 1 0 41888 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A1
timestamp 1669390400
transform -1 0 23296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__A2
timestamp 1669390400
transform 1 0 23520 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A1
timestamp 1669390400
transform 1 0 24640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A2
timestamp 1669390400
transform 1 0 23632 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A1
timestamp 1669390400
transform -1 0 11648 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__A2
timestamp 1669390400
transform -1 0 15120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A1
timestamp 1669390400
transform 1 0 25088 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__A2
timestamp 1669390400
transform 1 0 29008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__B1
timestamp 1669390400
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__B2
timestamp 1669390400
transform -1 0 34608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__B
timestamp 1669390400
transform -1 0 4032 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1669390400
transform -1 0 27888 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A2
timestamp 1669390400
transform 1 0 27216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A1
timestamp 1669390400
transform 1 0 25536 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A2
timestamp 1669390400
transform 1 0 25872 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__A1
timestamp 1669390400
transform 1 0 23072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__A2
timestamp 1669390400
transform 1 0 26096 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I0
timestamp 1669390400
transform 1 0 35952 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I1
timestamp 1669390400
transform 1 0 35056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I3
timestamp 1669390400
transform 1 0 36848 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__S0
timestamp 1669390400
transform 1 0 37296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__S1
timestamp 1669390400
transform 1 0 36400 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__I
timestamp 1669390400
transform -1 0 3360 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__A1
timestamp 1669390400
transform 1 0 28896 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__A2
timestamp 1669390400
transform -1 0 28672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A1
timestamp 1669390400
transform 1 0 28560 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A2
timestamp 1669390400
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A1
timestamp 1669390400
transform 1 0 31024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A2
timestamp 1669390400
transform 1 0 29792 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A1
timestamp 1669390400
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1669390400
transform 1 0 23632 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A2
timestamp 1669390400
transform 1 0 34384 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__B
timestamp 1669390400
transform 1 0 23184 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A1
timestamp 1669390400
transform -1 0 23856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A2
timestamp 1669390400
transform 1 0 23072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__B1
timestamp 1669390400
transform 1 0 20832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__B2
timestamp 1669390400
transform -1 0 24416 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A1
timestamp 1669390400
transform -1 0 26768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A2
timestamp 1669390400
transform 1 0 22624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A1
timestamp 1669390400
transform 1 0 32368 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A1
timestamp 1669390400
transform 1 0 30240 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A2
timestamp 1669390400
transform 1 0 32032 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A1
timestamp 1669390400
transform 1 0 37856 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A2
timestamp 1669390400
transform 1 0 38304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__B1
timestamp 1669390400
transform 1 0 36176 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__B2
timestamp 1669390400
transform -1 0 35728 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__C1
timestamp 1669390400
transform 1 0 35952 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__C2
timestamp 1669390400
transform -1 0 11984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A1
timestamp 1669390400
transform 1 0 4816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1669390400
transform -1 0 6832 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A1
timestamp 1669390400
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A2
timestamp 1669390400
transform 1 0 29568 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1669390400
transform 1 0 31920 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A2
timestamp 1669390400
transform 1 0 33040 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I0
timestamp 1669390400
transform 1 0 35952 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I1
timestamp 1669390400
transform -1 0 36064 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__I3
timestamp 1669390400
transform 1 0 36288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__S0
timestamp 1669390400
transform 1 0 37408 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__S1
timestamp 1669390400
transform 1 0 36736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1669390400
transform 1 0 35504 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A2
timestamp 1669390400
transform 1 0 35056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A1
timestamp 1669390400
transform 1 0 35056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A2
timestamp 1669390400
transform 1 0 34608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__B
timestamp 1669390400
transform 1 0 33488 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1669390400
transform 1 0 36512 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I0
timestamp 1669390400
transform 1 0 36736 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I1
timestamp 1669390400
transform -1 0 35728 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__I3
timestamp 1669390400
transform 1 0 37408 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__S0
timestamp 1669390400
transform 1 0 37856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__S1
timestamp 1669390400
transform -1 0 37184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1669390400
transform 1 0 37184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A2
timestamp 1669390400
transform 1 0 37856 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1669390400
transform -1 0 34160 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__A1
timestamp 1669390400
transform 1 0 34608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__A2
timestamp 1669390400
transform 1 0 32816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I0
timestamp 1669390400
transform 1 0 38080 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I1
timestamp 1669390400
transform -1 0 33264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__I3
timestamp 1669390400
transform 1 0 37632 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__S0
timestamp 1669390400
transform 1 0 38976 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__S1
timestamp 1669390400
transform 1 0 38528 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A1
timestamp 1669390400
transform 1 0 37408 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A2
timestamp 1669390400
transform 1 0 36400 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A1
timestamp 1669390400
transform 1 0 34160 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A1
timestamp 1669390400
transform 1 0 32816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A1
timestamp 1669390400
transform 1 0 34832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A2
timestamp 1669390400
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__B
timestamp 1669390400
transform 1 0 33936 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A1
timestamp 1669390400
transform 1 0 24080 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A2
timestamp 1669390400
transform 1 0 17136 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A1
timestamp 1669390400
transform 1 0 22176 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A2
timestamp 1669390400
transform 1 0 20720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__B1
timestamp 1669390400
transform 1 0 20272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__B2
timestamp 1669390400
transform 1 0 20160 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A1
timestamp 1669390400
transform 1 0 34384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A1
timestamp 1669390400
transform 1 0 2352 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A2
timestamp 1669390400
transform 1 0 11648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A1
timestamp 1669390400
transform -1 0 2464 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__A2
timestamp 1669390400
transform 1 0 2688 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__B
timestamp 1669390400
transform 1 0 3136 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A1
timestamp 1669390400
transform -1 0 8736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A2
timestamp 1669390400
transform -1 0 2912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A1
timestamp 1669390400
transform -1 0 12544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A2
timestamp 1669390400
transform -1 0 4704 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A1
timestamp 1669390400
transform -1 0 16016 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A2
timestamp 1669390400
transform 1 0 6272 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__B2
timestamp 1669390400
transform -1 0 15568 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1669390400
transform 1 0 20832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A2
timestamp 1669390400
transform -1 0 20496 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__A1
timestamp 1669390400
transform -1 0 3808 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__A2
timestamp 1669390400
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__C
timestamp 1669390400
transform -1 0 4704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A1
timestamp 1669390400
transform 1 0 4816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A2
timestamp 1669390400
transform 1 0 8064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A3
timestamp 1669390400
transform 1 0 4032 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A1
timestamp 1669390400
transform -1 0 4480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A2
timestamp 1669390400
transform 1 0 3808 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__B1
timestamp 1669390400
transform -1 0 4256 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__B2
timestamp 1669390400
transform -1 0 3136 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__C1
timestamp 1669390400
transform 1 0 3360 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__C2
timestamp 1669390400
transform 1 0 4704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A1
timestamp 1669390400
transform -1 0 6384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A2
timestamp 1669390400
transform -1 0 6048 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A1
timestamp 1669390400
transform 1 0 8960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A2
timestamp 1669390400
transform 1 0 8512 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1669390400
transform -1 0 2016 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A2
timestamp 1669390400
transform 1 0 3136 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A2
timestamp 1669390400
transform -1 0 2352 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A1
timestamp 1669390400
transform -1 0 8288 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A2
timestamp 1669390400
transform -1 0 6944 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A1
timestamp 1669390400
transform -1 0 7840 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A2
timestamp 1669390400
transform 1 0 4480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A1
timestamp 1669390400
transform -1 0 7952 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__CLK
timestamp 1669390400
transform 1 0 41328 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__D
timestamp 1669390400
transform 1 0 40880 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__CLK
timestamp 1669390400
transform -1 0 37072 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__D
timestamp 1669390400
transform 1 0 35280 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__CLK
timestamp 1669390400
transform -1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__D
timestamp 1669390400
transform -1 0 5152 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__CLK
timestamp 1669390400
transform 1 0 39200 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__D
timestamp 1669390400
transform 1 0 38752 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__CLK
timestamp 1669390400
transform 1 0 38752 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__D
timestamp 1669390400
transform -1 0 9632 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__CLK
timestamp 1669390400
transform -1 0 25984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__D
timestamp 1669390400
transform -1 0 9856 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__CLK
timestamp 1669390400
transform -1 0 2016 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__D
timestamp 1669390400
transform -1 0 2240 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__CLK
timestamp 1669390400
transform 1 0 18928 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__D
timestamp 1669390400
transform -1 0 18256 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__CLK
timestamp 1669390400
transform 1 0 5376 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__CLK
timestamp 1669390400
transform 1 0 15344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__D
timestamp 1669390400
transform -1 0 2016 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__CLK
timestamp 1669390400
transform 1 0 38640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__D
timestamp 1669390400
transform 1 0 38192 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__CLK
timestamp 1669390400
transform 1 0 13328 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__D
timestamp 1669390400
transform -1 0 2464 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__CLK
timestamp 1669390400
transform 1 0 39648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__D
timestamp 1669390400
transform -1 0 3696 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__CLK
timestamp 1669390400
transform 1 0 15120 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__D
timestamp 1669390400
transform -1 0 9856 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__CLK
timestamp 1669390400
transform 1 0 25312 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__D
timestamp 1669390400
transform -1 0 25088 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__CLK
timestamp 1669390400
transform -1 0 7280 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__D
timestamp 1669390400
transform 1 0 4928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__CLK
timestamp 1669390400
transform -1 0 10304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__D
timestamp 1669390400
transform -1 0 9408 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__CLK
timestamp 1669390400
transform 1 0 35728 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__D
timestamp 1669390400
transform -1 0 22064 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__CLK
timestamp 1669390400
transform 1 0 3136 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__CLK
timestamp 1669390400
transform 1 0 38304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__D
timestamp 1669390400
transform 1 0 37856 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__CLK
timestamp 1669390400
transform 1 0 40992 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__D
timestamp 1669390400
transform -1 0 2576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__CLK
timestamp 1669390400
transform 1 0 4480 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__D
timestamp 1669390400
transform -1 0 2464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__CLK
timestamp 1669390400
transform 1 0 21280 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__D
timestamp 1669390400
transform -1 0 21952 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__CLK
timestamp 1669390400
transform 1 0 37296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__CLK
timestamp 1669390400
transform 1 0 39648 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__CLK
timestamp 1669390400
transform 1 0 22624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__CLK
timestamp 1669390400
transform 1 0 9408 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__D
timestamp 1669390400
transform -1 0 8736 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__CLK
timestamp 1669390400
transform 1 0 14672 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__D
timestamp 1669390400
transform 1 0 40768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__CLK
timestamp 1669390400
transform 1 0 40320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__CLK
timestamp 1669390400
transform 1 0 14000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__D
timestamp 1669390400
transform -1 0 2912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__CLK
timestamp 1669390400
transform -1 0 11760 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__D
timestamp 1669390400
transform -1 0 10528 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__CLK
timestamp 1669390400
transform 1 0 40096 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__542__D
timestamp 1669390400
transform 1 0 41440 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__CLK
timestamp 1669390400
transform 1 0 7280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__D
timestamp 1669390400
transform -1 0 4480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__CLK
timestamp 1669390400
transform 1 0 39536 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__D
timestamp 1669390400
transform -1 0 2912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__CLK
timestamp 1669390400
transform 1 0 14000 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__CLK
timestamp 1669390400
transform -1 0 2016 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__D
timestamp 1669390400
transform -1 0 9856 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__CLK
timestamp 1669390400
transform 1 0 23520 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__D
timestamp 1669390400
transform -1 0 19264 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__CLK
timestamp 1669390400
transform 1 0 40544 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__D
timestamp 1669390400
transform 1 0 40096 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform -1 0 2240 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 4032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 52640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 55104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 60032 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 63952 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 67872 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 72576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform 1 0 16240 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform -1 0 2128 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 3024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 38304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 39200 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 35952 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 37632 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 42000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform 1 0 48720 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform 1 0 77168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 74368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1669390400
transform -1 0 4368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output25_I
timestamp 1669390400
transform -1 0 72688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2240 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23
timestamp 1669390400
transform 1 0 3920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45
timestamp 1669390400
transform 1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49
timestamp 1669390400
transform 1 0 6832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65
timestamp 1669390400
transform 1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1669390400
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_123
timestamp 1669390400
transform 1 0 15120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127
timestamp 1669390400
transform 1 0 15568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_129
timestamp 1669390400
transform 1 0 15792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_132
timestamp 1669390400
transform 1 0 16128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_157
timestamp 1669390400
transform 1 0 18928 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1669390400
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_192
timestamp 1669390400
transform 1 0 22848 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_208
timestamp 1669390400
transform 1 0 24640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_216
timestamp 1669390400
transform 1 0 25536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_218
timestamp 1669390400
transform 1 0 25760 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_233
timestamp 1669390400
transform 1 0 27440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_241
timestamp 1669390400
transform 1 0 28336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_255
timestamp 1669390400
transform 1 0 29904 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_259
timestamp 1669390400
transform 1 0 30352 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_275
timestamp 1669390400
transform 1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1669390400
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_367
timestamp 1669390400
transform 1 0 42448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_383
timestamp 1669390400
transform 1 0 44240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_402
timestamp 1669390400
transform 1 0 46368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_426
timestamp 1669390400
transform 1 0 49056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_428
timestamp 1669390400
transform 1 0 49280 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_443
timestamp 1669390400
transform 1 0 50960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_447
timestamp 1669390400
transform 1 0 51408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_450
timestamp 1669390400
transform 1 0 51744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_466
timestamp 1669390400
transform 1 0 53536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_470
timestamp 1669390400
transform 1 0 53984 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_485
timestamp 1669390400
transform 1 0 55664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1669390400
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_577
timestamp 1669390400
transform 1 0 65968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_593
timestamp 1669390400
transform 1 0 67760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_612
timestamp 1669390400
transform 1 0 69888 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_628
timestamp 1669390400
transform 1 0 71680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_634
timestamp 1669390400
transform 1 0 72352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_637
timestamp 1669390400
transform 1 0 72688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_653
timestamp 1669390400
transform 1 0 74480 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_661
timestamp 1669390400
transform 1 0 75376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_683
timestamp 1669390400
transform 1 0 77840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_687
timestamp 1669390400
transform 1 0 78288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_34
timestamp 1669390400
transform 1 0 5152 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_50
timestamp 1669390400
transform 1 0 6944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_58
timestamp 1669390400
transform 1 0 7840 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_81
timestamp 1669390400
transform 1 0 10416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_85
timestamp 1669390400
transform 1 0 10864 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_87
timestamp 1669390400
transform 1 0 11088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_96
timestamp 1669390400
transform 1 0 12096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_100
timestamp 1669390400
transform 1 0 12544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_112
timestamp 1669390400
transform 1 0 13888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_116
timestamp 1669390400
transform 1 0 14336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_120
timestamp 1669390400
transform 1 0 14784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_130
timestamp 1669390400
transform 1 0 15904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_138
timestamp 1669390400
transform 1 0 16800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_160
timestamp 1669390400
transform 1 0 19264 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_168
timestamp 1669390400
transform 1 0 20160 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_200
timestamp 1669390400
transform 1 0 23744 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_223
timestamp 1669390400
transform 1 0 26320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_229
timestamp 1669390400
transform 1 0 26992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_233
timestamp 1669390400
transform 1 0 27440 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_243
timestamp 1669390400
transform 1 0 28560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_247
timestamp 1669390400
transform 1 0 29008 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_254
timestamp 1669390400
transform 1 0 29792 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_270
timestamp 1669390400
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_278
timestamp 1669390400
transform 1 0 32480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_282
timestamp 1669390400
transform 1 0 32928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_290
timestamp 1669390400
transform 1 0 33824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_292
timestamp 1669390400
transform 1 0 34048 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_299
timestamp 1669390400
transform 1 0 34832 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_315
timestamp 1669390400
transform 1 0 36624 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_323
timestamp 1669390400
transform 1 0 37520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_327
timestamp 1669390400
transform 1 0 37968 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_335
timestamp 1669390400
transform 1 0 38864 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_351
timestamp 1669390400
transform 1 0 40656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_373
timestamp 1669390400
transform 1 0 43120 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_381
timestamp 1669390400
transform 1 0 44016 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_413
timestamp 1669390400
transform 1 0 47600 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_435
timestamp 1669390400
transform 1 0 50064 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_439
timestamp 1669390400
transform 1 0 50512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_443
timestamp 1669390400
transform 1 0 50960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_447
timestamp 1669390400
transform 1 0 51408 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_457
timestamp 1669390400
transform 1 0 52528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_467
timestamp 1669390400
transform 1 0 53648 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_475
timestamp 1669390400
transform 1 0 54544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_483
timestamp 1669390400
transform 1 0 55440 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_491
timestamp 1669390400
transform 1 0 56336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1669390400
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_503
timestamp 1669390400
transform 1 0 57680 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_510
timestamp 1669390400
transform 1 0 58464 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_542
timestamp 1669390400
transform 1 0 62048 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_558
timestamp 1669390400
transform 1 0 63840 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_566
timestamp 1669390400
transform 1 0 64736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_573
timestamp 1669390400
transform 1 0 65520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_581
timestamp 1669390400
transform 1 0 66416 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_613
timestamp 1669390400
transform 1 0 70000 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_629
timestamp 1669390400
transform 1 0 71792 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_637
timestamp 1669390400
transform 1 0 72688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_649
timestamp 1669390400
transform 1 0 74032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_651
timestamp 1669390400
transform 1 0 74256 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_654
timestamp 1669390400
transform 1 0 74592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_670
timestamp 1669390400
transform 1 0 76384 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_686
timestamp 1669390400
transform 1 0 78176 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_69
timestamp 1669390400
transform 1 0 9072 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_85
timestamp 1669390400
transform 1 0 10864 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_87
timestamp 1669390400
transform 1 0 11088 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_94
timestamp 1669390400
transform 1 0 11872 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_102
timestamp 1669390400
transform 1 0 12768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_183
timestamp 1669390400
transform 1 0 21840 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_185
timestamp 1669390400
transform 1 0 22064 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_188
timestamp 1669390400
transform 1 0 22400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_192
timestamp 1669390400
transform 1 0 22848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_202
timestamp 1669390400
transform 1 0 23968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_210
timestamp 1669390400
transform 1 0 24864 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_242
timestamp 1669390400
transform 1 0 28448 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_246
timestamp 1669390400
transform 1 0 28896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_266
timestamp 1669390400
transform 1 0 31136 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_276
timestamp 1669390400
transform 1 0 32256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_280
timestamp 1669390400
transform 1 0 32704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_290
timestamp 1669390400
transform 1 0 33824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_292
timestamp 1669390400
transform 1 0 34048 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_295
timestamp 1669390400
transform 1 0 34384 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_305
timestamp 1669390400
transform 1 0 35504 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_313
timestamp 1669390400
transform 1 0 36400 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_317
timestamp 1669390400
transform 1 0 36848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_337
timestamp 1669390400
transform 1 0 39088 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_339
timestamp 1669390400
transform 1 0 39312 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_342
timestamp 1669390400
transform 1 0 39648 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_346
timestamp 1669390400
transform 1 0 40096 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_356
timestamp 1669390400
transform 1 0 41216 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1669390400
transform 1 0 44800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_400
timestamp 1669390400
transform 1 0 46144 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_404
timestamp 1669390400
transform 1 0 46592 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_407
timestamp 1669390400
transform 1 0 46928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_411
timestamp 1669390400
transform 1 0 47376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_421
timestamp 1669390400
transform 1 0 48496 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_453
timestamp 1669390400
transform 1 0 52080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_457
timestamp 1669390400
transform 1 0 52528 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_466
timestamp 1669390400
transform 1 0 53536 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_530
timestamp 1669390400
transform 1 0 60704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_598
timestamp 1669390400
transform 1 0 68320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_669
timestamp 1669390400
transform 1 0 76272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1669390400
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_684
timestamp 1669390400
transform 1 0 77952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_81
timestamp 1669390400
transform 1 0 10416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_93
timestamp 1669390400
transform 1 0 11760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_97
timestamp 1669390400
transform 1 0 12208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_101
timestamp 1669390400
transform 1 0 12656 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_109
timestamp 1669390400
transform 1 0 13552 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_113
timestamp 1669390400
transform 1 0 14000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_117
timestamp 1669390400
transform 1 0 14448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_127
timestamp 1669390400
transform 1 0 15568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_135
timestamp 1669390400
transform 1 0 16464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_139
timestamp 1669390400
transform 1 0 16912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_148
timestamp 1669390400
transform 1 0 17920 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_151
timestamp 1669390400
transform 1 0 18256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_161
timestamp 1669390400
transform 1 0 19376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_165
timestamp 1669390400
transform 1 0 19824 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_197
timestamp 1669390400
transform 1 0 23408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_290
timestamp 1669390400
transform 1 0 33824 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_292
timestamp 1669390400
transform 1 0 34048 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_295
timestamp 1669390400
transform 1 0 34384 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_327
timestamp 1669390400
transform 1 0 37968 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_343
timestamp 1669390400
transform 1 0 39760 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_351
timestamp 1669390400
transform 1 0 40656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_444
timestamp 1669390400
transform 1 0 51072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_447
timestamp 1669390400
transform 1 0 51408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_451
timestamp 1669390400
transform 1 0 51856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_461
timestamp 1669390400
transform 1 0 52976 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_493
timestamp 1669390400
transform 1 0 56560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_673
timestamp 1669390400
transform 1 0 76720 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_681
timestamp 1669390400
transform 1 0 77616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_685
timestamp 1669390400
transform 1 0 78064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_687
timestamp 1669390400
transform 1 0 78288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1669390400
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_684
timestamp 1669390400
transform 1 0 77952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_673
timestamp 1669390400
transform 1 0 76720 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_681
timestamp 1669390400
transform 1 0 77616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_685
timestamp 1669390400
transform 1 0 78064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_687
timestamp 1669390400
transform 1 0 78288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_684
timestamp 1669390400
transform 1 0 77952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_673
timestamp 1669390400
transform 1 0 76720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_681
timestamp 1669390400
transform 1 0 77616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_685
timestamp 1669390400
transform 1 0 78064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_687
timestamp 1669390400
transform 1 0 78288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_684
timestamp 1669390400
transform 1 0 77952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_673
timestamp 1669390400
transform 1 0 76720 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_681
timestamp 1669390400
transform 1 0 77616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_685
timestamp 1669390400
transform 1 0 78064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_687
timestamp 1669390400
transform 1 0 78288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_684
timestamp 1669390400
transform 1 0 77952 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_673
timestamp 1669390400
transform 1 0 76720 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_681
timestamp 1669390400
transform 1 0 77616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_685
timestamp 1669390400
transform 1 0 78064 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_687
timestamp 1669390400
transform 1 0 78288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_684
timestamp 1669390400
transform 1 0 77952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_673
timestamp 1669390400
transform 1 0 76720 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_681
timestamp 1669390400
transform 1 0 77616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_685
timestamp 1669390400
transform 1 0 78064 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_687
timestamp 1669390400
transform 1 0 78288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_684
timestamp 1669390400
transform 1 0 77952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_673
timestamp 1669390400
transform 1 0 76720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_681
timestamp 1669390400
transform 1 0 77616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_685
timestamp 1669390400
transform 1 0 78064 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_687
timestamp 1669390400
transform 1 0 78288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_684
timestamp 1669390400
transform 1 0 77952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_673
timestamp 1669390400
transform 1 0 76720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_681
timestamp 1669390400
transform 1 0 77616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_685
timestamp 1669390400
transform 1 0 78064 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_687
timestamp 1669390400
transform 1 0 78288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_684
timestamp 1669390400
transform 1 0 77952 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_673
timestamp 1669390400
transform 1 0 76720 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_681
timestamp 1669390400
transform 1 0 77616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_685
timestamp 1669390400
transform 1 0 78064 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_687
timestamp 1669390400
transform 1 0 78288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_684
timestamp 1669390400
transform 1 0 77952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_673
timestamp 1669390400
transform 1 0 76720 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_681
timestamp 1669390400
transform 1 0 77616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_685
timestamp 1669390400
transform 1 0 78064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_687
timestamp 1669390400
transform 1 0 78288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_684
timestamp 1669390400
transform 1 0 77952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_673
timestamp 1669390400
transform 1 0 76720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_681
timestamp 1669390400
transform 1 0 77616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_685
timestamp 1669390400
transform 1 0 78064 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1669390400
transform 1 0 78288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_684
timestamp 1669390400
transform 1 0 77952 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_673
timestamp 1669390400
transform 1 0 76720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_681
timestamp 1669390400
transform 1 0 77616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_685
timestamp 1669390400
transform 1 0 78064 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1669390400
transform 1 0 78288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_684
timestamp 1669390400
transform 1 0 77952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_673
timestamp 1669390400
transform 1 0 76720 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_681
timestamp 1669390400
transform 1 0 77616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_685
timestamp 1669390400
transform 1 0 78064 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1669390400
transform 1 0 78288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_684
timestamp 1669390400
transform 1 0 77952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_673
timestamp 1669390400
transform 1 0 76720 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_681
timestamp 1669390400
transform 1 0 77616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_685
timestamp 1669390400
transform 1 0 78064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1669390400
transform 1 0 78288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_684
timestamp 1669390400
transform 1 0 77952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_673
timestamp 1669390400
transform 1 0 76720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_681
timestamp 1669390400
transform 1 0 77616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_685
timestamp 1669390400
transform 1 0 78064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1669390400
transform 1 0 78288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_684
timestamp 1669390400
transform 1 0 77952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_673
timestamp 1669390400
transform 1 0 76720 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_681
timestamp 1669390400
transform 1 0 77616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_685
timestamp 1669390400
transform 1 0 78064 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1669390400
transform 1 0 78288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_684
timestamp 1669390400
transform 1 0 77952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_673
timestamp 1669390400
transform 1 0 76720 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_681
timestamp 1669390400
transform 1 0 77616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_685
timestamp 1669390400
transform 1 0 78064 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1669390400
transform 1 0 78288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1669390400
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_684
timestamp 1669390400
transform 1 0 77952 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1669390400
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1669390400
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_673
timestamp 1669390400
transform 1 0 76720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_681
timestamp 1669390400
transform 1 0 77616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_685
timestamp 1669390400
transform 1 0 78064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1669390400
transform 1 0 78288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1669390400
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1669390400
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_684
timestamp 1669390400
transform 1 0 77952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1669390400
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1669390400
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_673
timestamp 1669390400
transform 1 0 76720 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_681
timestamp 1669390400
transform 1 0 77616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_685
timestamp 1669390400
transform 1 0 78064 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1669390400
transform 1 0 78288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1669390400
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1669390400
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1669390400
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1669390400
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_684
timestamp 1669390400
transform 1 0 77952 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1669390400
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1669390400
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_673
timestamp 1669390400
transform 1 0 76720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_681
timestamp 1669390400
transform 1 0 77616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_685
timestamp 1669390400
transform 1 0 78064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1669390400
transform 1 0 78288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_124
timestamp 1669390400
transform 1 0 15232 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_132
timestamp 1669390400
transform 1 0 16128 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_136
timestamp 1669390400
transform 1 0 16576 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_138
timestamp 1669390400
transform 1 0 16800 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_141
timestamp 1669390400
transform 1 0 17136 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_149
timestamp 1669390400
transform 1 0 18032 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_165
timestamp 1669390400
transform 1 0 19824 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_173
timestamp 1669390400
transform 1 0 20720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1669390400
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1669390400
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1669390400
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1669390400
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_669
timestamp 1669390400
transform 1 0 76272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1669390400
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_676
timestamp 1669390400
transform 1 0 77056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_684
timestamp 1669390400
transform 1 0 77952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_563
timestamp 1669390400
transform 1 0 64400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1669390400
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1669390400
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1669390400
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1669390400
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_641
timestamp 1669390400
transform 1 0 73136 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_673
timestamp 1669390400
transform 1 0 76720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_681
timestamp 1669390400
transform 1 0 77616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_685
timestamp 1669390400
transform 1 0 78064 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_687
timestamp 1669390400
transform 1 0 78288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_527
timestamp 1669390400
transform 1 0 60368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1669390400
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_598
timestamp 1669390400
transform 1 0 68320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1669390400
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1669390400
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_669
timestamp 1669390400
transform 1 0 76272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1669390400
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_676
timestamp 1669390400
transform 1 0 77056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_684
timestamp 1669390400
transform 1 0 77952 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1669390400
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_563
timestamp 1669390400
transform 1 0 64400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1669390400
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1669390400
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1669390400
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1669390400
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_641
timestamp 1669390400
transform 1 0 73136 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_673
timestamp 1669390400
transform 1 0 76720 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_681
timestamp 1669390400
transform 1 0 77616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_685
timestamp 1669390400
transform 1 0 78064 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_687
timestamp 1669390400
transform 1 0 78288 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1669390400
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_527
timestamp 1669390400
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1669390400
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1669390400
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1669390400
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_605
timestamp 1669390400
transform 1 0 69104 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_669
timestamp 1669390400
transform 1 0 76272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1669390400
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_676
timestamp 1669390400
transform 1 0 77056 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_684
timestamp 1669390400
transform 1 0 77952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_421
timestamp 1669390400
transform 1 0 48496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1669390400
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1669390400
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1669390400
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1669390400
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1669390400
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_641
timestamp 1669390400
transform 1 0 73136 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_673
timestamp 1669390400
transform 1 0 76720 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_681
timestamp 1669390400
transform 1 0 77616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_685
timestamp 1669390400
transform 1 0 78064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_687
timestamp 1669390400
transform 1 0 78288 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_527
timestamp 1669390400
transform 1 0 60368 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1669390400
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_598
timestamp 1669390400
transform 1 0 68320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1669390400
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1669390400
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_669
timestamp 1669390400
transform 1 0 76272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1669390400
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_676
timestamp 1669390400
transform 1 0 77056 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_684
timestamp 1669390400
transform 1 0 77952 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1669390400
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1669390400
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_563
timestamp 1669390400
transform 1 0 64400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1669390400
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1669390400
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1669390400
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1669390400
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_641
timestamp 1669390400
transform 1 0 73136 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_673
timestamp 1669390400
transform 1 0 76720 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_681
timestamp 1669390400
transform 1 0 77616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_685
timestamp 1669390400
transform 1 0 78064 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_687
timestamp 1669390400
transform 1 0 78288 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1669390400
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_527
timestamp 1669390400
transform 1 0 60368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1669390400
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_598
timestamp 1669390400
transform 1 0 68320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1669390400
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1669390400
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_669
timestamp 1669390400
transform 1 0 76272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1669390400
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_676
timestamp 1669390400
transform 1 0 77056 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_684
timestamp 1669390400
transform 1 0 77952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_421
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_563
timestamp 1669390400
transform 1 0 64400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1669390400
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1669390400
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_634
timestamp 1669390400
transform 1 0 72352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1669390400
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_641
timestamp 1669390400
transform 1 0 73136 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_673
timestamp 1669390400
transform 1 0 76720 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_681
timestamp 1669390400
transform 1 0 77616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_685
timestamp 1669390400
transform 1 0 78064 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_687
timestamp 1669390400
transform 1 0 78288 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_456
timestamp 1669390400
transform 1 0 52416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1669390400
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1669390400
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_598
timestamp 1669390400
transform 1 0 68320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1669390400
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1669390400
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_669
timestamp 1669390400
transform 1 0 76272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1669390400
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_676
timestamp 1669390400
transform 1 0 77056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_684
timestamp 1669390400
transform 1 0 77952 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_563
timestamp 1669390400
transform 1 0 64400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1669390400
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1669390400
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_634
timestamp 1669390400
transform 1 0 72352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1669390400
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_641
timestamp 1669390400
transform 1 0 73136 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_673
timestamp 1669390400
transform 1 0 76720 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_681
timestamp 1669390400
transform 1 0 77616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_685
timestamp 1669390400
transform 1 0 78064 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_687
timestamp 1669390400
transform 1 0 78288 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_527
timestamp 1669390400
transform 1 0 60368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1669390400
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_598
timestamp 1669390400
transform 1 0 68320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1669390400
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_605
timestamp 1669390400
transform 1 0 69104 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_669
timestamp 1669390400
transform 1 0 76272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1669390400
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_676
timestamp 1669390400
transform 1 0 77056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_684
timestamp 1669390400
transform 1 0 77952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_563
timestamp 1669390400
transform 1 0 64400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1669390400
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1669390400
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_634
timestamp 1669390400
transform 1 0 72352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1669390400
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_641
timestamp 1669390400
transform 1 0 73136 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_673
timestamp 1669390400
transform 1 0 76720 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_681
timestamp 1669390400
transform 1 0 77616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_685
timestamp 1669390400
transform 1 0 78064 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_687
timestamp 1669390400
transform 1 0 78288 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_527
timestamp 1669390400
transform 1 0 60368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1669390400
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_598
timestamp 1669390400
transform 1 0 68320 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1669390400
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_605
timestamp 1669390400
transform 1 0 69104 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_669
timestamp 1669390400
transform 1 0 76272 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1669390400
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_676
timestamp 1669390400
transform 1 0 77056 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_684
timestamp 1669390400
transform 1 0 77952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_421
timestamp 1669390400
transform 1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_563
timestamp 1669390400
transform 1 0 64400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1669390400
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_570
timestamp 1669390400
transform 1 0 65184 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_634
timestamp 1669390400
transform 1 0 72352 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1669390400
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_641
timestamp 1669390400
transform 1 0 73136 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_673
timestamp 1669390400
transform 1 0 76720 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_681
timestamp 1669390400
transform 1 0 77616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_685
timestamp 1669390400
transform 1 0 78064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_687
timestamp 1669390400
transform 1 0 78288 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_456
timestamp 1669390400
transform 1 0 52416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_527
timestamp 1669390400
transform 1 0 60368 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1669390400
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_598
timestamp 1669390400
transform 1 0 68320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1669390400
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_605
timestamp 1669390400
transform 1 0 69104 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_669
timestamp 1669390400
transform 1 0 76272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_673
timestamp 1669390400
transform 1 0 76720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_676
timestamp 1669390400
transform 1 0 77056 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_684
timestamp 1669390400
transform 1 0 77952 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1669390400
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_563
timestamp 1669390400
transform 1 0 64400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1669390400
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_570
timestamp 1669390400
transform 1 0 65184 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_634
timestamp 1669390400
transform 1 0 72352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1669390400
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_641
timestamp 1669390400
transform 1 0 73136 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_673
timestamp 1669390400
transform 1 0 76720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_681
timestamp 1669390400
transform 1 0 77616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_685
timestamp 1669390400
transform 1 0 78064 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_687
timestamp 1669390400
transform 1 0 78288 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1669390400
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_527
timestamp 1669390400
transform 1 0 60368 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1669390400
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_598
timestamp 1669390400
transform 1 0 68320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1669390400
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_605
timestamp 1669390400
transform 1 0 69104 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_669
timestamp 1669390400
transform 1 0 76272 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_673
timestamp 1669390400
transform 1 0 76720 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_676
timestamp 1669390400
transform 1 0 77056 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_684
timestamp 1669390400
transform 1 0 77952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1669390400
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_492
timestamp 1669390400
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_563
timestamp 1669390400
transform 1 0 64400 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_567
timestamp 1669390400
transform 1 0 64848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1669390400
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_634
timestamp 1669390400
transform 1 0 72352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1669390400
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_641
timestamp 1669390400
transform 1 0 73136 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_673
timestamp 1669390400
transform 1 0 76720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_681
timestamp 1669390400
transform 1 0 77616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_685
timestamp 1669390400
transform 1 0 78064 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_687
timestamp 1669390400
transform 1 0 78288 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_456
timestamp 1669390400
transform 1 0 52416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_527
timestamp 1669390400
transform 1 0 60368 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1669390400
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_598
timestamp 1669390400
transform 1 0 68320 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_602
timestamp 1669390400
transform 1 0 68768 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_605
timestamp 1669390400
transform 1 0 69104 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_669
timestamp 1669390400
transform 1 0 76272 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1669390400
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_676
timestamp 1669390400
transform 1 0 77056 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_684
timestamp 1669390400
transform 1 0 77952 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1669390400
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_563
timestamp 1669390400
transform 1 0 64400 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1669390400
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1669390400
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_634
timestamp 1669390400
transform 1 0 72352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1669390400
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_641
timestamp 1669390400
transform 1 0 73136 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_673
timestamp 1669390400
transform 1 0 76720 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_681
timestamp 1669390400
transform 1 0 77616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_685
timestamp 1669390400
transform 1 0 78064 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_687
timestamp 1669390400
transform 1 0 78288 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_527
timestamp 1669390400
transform 1 0 60368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_531
timestamp 1669390400
transform 1 0 60816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_598
timestamp 1669390400
transform 1 0 68320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1669390400
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_605
timestamp 1669390400
transform 1 0 69104 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_669
timestamp 1669390400
transform 1 0 76272 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1669390400
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_676
timestamp 1669390400
transform 1 0 77056 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_684
timestamp 1669390400
transform 1 0 77952 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_563
timestamp 1669390400
transform 1 0 64400 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_567
timestamp 1669390400
transform 1 0 64848 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1669390400
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_634
timestamp 1669390400
transform 1 0 72352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1669390400
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_641
timestamp 1669390400
transform 1 0 73136 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_673
timestamp 1669390400
transform 1 0 76720 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_681
timestamp 1669390400
transform 1 0 77616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_685
timestamp 1669390400
transform 1 0 78064 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_687
timestamp 1669390400
transform 1 0 78288 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_257
timestamp 1669390400
transform 1 0 30128 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_289
timestamp 1669390400
transform 1 0 33712 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_305
timestamp 1669390400
transform 1 0 35504 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_313
timestamp 1669390400
transform 1 0 36400 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_317
timestamp 1669390400
transform 1 0 36848 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_456
timestamp 1669390400
transform 1 0 52416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_527
timestamp 1669390400
transform 1 0 60368 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1669390400
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_598
timestamp 1669390400
transform 1 0 68320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1669390400
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_605
timestamp 1669390400
transform 1 0 69104 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_669
timestamp 1669390400
transform 1 0 76272 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1669390400
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_676
timestamp 1669390400
transform 1 0 77056 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_684
timestamp 1669390400
transform 1 0 77952 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1669390400
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1669390400
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1669390400
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_563
timestamp 1669390400
transform 1 0 64400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_567
timestamp 1669390400
transform 1 0 64848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1669390400
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_634
timestamp 1669390400
transform 1 0 72352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1669390400
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_641
timestamp 1669390400
transform 1 0 73136 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_673
timestamp 1669390400
transform 1 0 76720 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_681
timestamp 1669390400
transform 1 0 77616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_685
timestamp 1669390400
transform 1 0 78064 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_687
timestamp 1669390400
transform 1 0 78288 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1669390400
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_69
timestamp 1669390400
transform 1 0 9072 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_72
timestamp 1669390400
transform 1 0 9408 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_76
timestamp 1669390400
transform 1 0 9856 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_80
timestamp 1669390400
transform 1 0 10304 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_96
timestamp 1669390400
transform 1 0 12096 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_98
timestamp 1669390400
transform 1 0 12320 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_101
timestamp 1669390400
transform 1 0 12656 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_111
timestamp 1669390400
transform 1 0 13776 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_115
timestamp 1669390400
transform 1 0 14224 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_147
timestamp 1669390400
transform 1 0 17808 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_163
timestamp 1669390400
transform 1 0 19600 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_171
timestamp 1669390400
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_175
timestamp 1669390400
transform 1 0 20944 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1669390400
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1669390400
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1669390400
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1669390400
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_456
timestamp 1669390400
transform 1 0 52416 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_527
timestamp 1669390400
transform 1 0 60368 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_531
timestamp 1669390400
transform 1 0 60816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_598
timestamp 1669390400
transform 1 0 68320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1669390400
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_605
timestamp 1669390400
transform 1 0 69104 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_669
timestamp 1669390400
transform 1 0 76272 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_673
timestamp 1669390400
transform 1 0 76720 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_676
timestamp 1669390400
transform 1 0 77056 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_684
timestamp 1669390400
transform 1 0 77952 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_34
timestamp 1669390400
transform 1 0 5152 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_50
timestamp 1669390400
transform 1 0 6944 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_52
timestamp 1669390400
transform 1 0 7168 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_55
timestamp 1669390400
transform 1 0 7504 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_59
timestamp 1669390400
transform 1 0 7952 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_63
timestamp 1669390400
transform 1 0 8400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_69
timestamp 1669390400
transform 1 0 9072 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_76
timestamp 1669390400
transform 1 0 9856 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_82
timestamp 1669390400
transform 1 0 10528 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_88
timestamp 1669390400
transform 1 0 11200 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_92
timestamp 1669390400
transform 1 0 11648 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_96
timestamp 1669390400
transform 1 0 12096 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_100
timestamp 1669390400
transform 1 0 12544 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_102
timestamp 1669390400
transform 1 0 12768 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_105
timestamp 1669390400
transform 1 0 13104 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_109
timestamp 1669390400
transform 1 0 13552 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_113
timestamp 1669390400
transform 1 0 14000 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_117
timestamp 1669390400
transform 1 0 14448 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_121
timestamp 1669390400
transform 1 0 14896 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_125
timestamp 1669390400
transform 1 0 15344 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1669390400
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1669390400
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1669390400
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1669390400
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1669390400
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1669390400
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1669390400
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_492
timestamp 1669390400
transform 1 0 56448 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1669390400
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_563
timestamp 1669390400
transform 1 0 64400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1669390400
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1669390400
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_634
timestamp 1669390400
transform 1 0 72352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1669390400
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_641
timestamp 1669390400
transform 1 0 73136 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_673
timestamp 1669390400
transform 1 0 76720 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_681
timestamp 1669390400
transform 1 0 77616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_685
timestamp 1669390400
transform 1 0 78064 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_687
timestamp 1669390400
transform 1 0 78288 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_18
timestamp 1669390400
transform 1 0 3360 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_22
timestamp 1669390400
transform 1 0 3808 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_25
timestamp 1669390400
transform 1 0 4144 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_33
timestamp 1669390400
transform 1 0 5040 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_41
timestamp 1669390400
transform 1 0 5936 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_45
timestamp 1669390400
transform 1 0 6384 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_49
timestamp 1669390400
transform 1 0 6832 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_51
timestamp 1669390400
transform 1 0 7056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_54
timestamp 1669390400
transform 1 0 7392 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_58
timestamp 1669390400
transform 1 0 7840 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_62
timestamp 1669390400
transform 1 0 8288 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_68
timestamp 1669390400
transform 1 0 8960 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_72
timestamp 1669390400
transform 1 0 9408 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_76
timestamp 1669390400
transform 1 0 9856 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_80
timestamp 1669390400
transform 1 0 10304 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_84
timestamp 1669390400
transform 1 0 10752 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_86
timestamp 1669390400
transform 1 0 10976 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_89
timestamp 1669390400
transform 1 0 11312 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_93
timestamp 1669390400
transform 1 0 11760 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_97
timestamp 1669390400
transform 1 0 12208 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_101
timestamp 1669390400
transform 1 0 12656 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_111
timestamp 1669390400
transform 1 0 13776 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_115
timestamp 1669390400
transform 1 0 14224 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_119
timestamp 1669390400
transform 1 0 14672 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_123
timestamp 1669390400
transform 1 0 15120 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_127
timestamp 1669390400
transform 1 0 15568 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_131
timestamp 1669390400
transform 1 0 16016 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_135
timestamp 1669390400
transform 1 0 16464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_139
timestamp 1669390400
transform 1 0 16912 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_143
timestamp 1669390400
transform 1 0 17360 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_147
timestamp 1669390400
transform 1 0 17808 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_151
timestamp 1669390400
transform 1 0 18256 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_159
timestamp 1669390400
transform 1 0 19152 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_165
timestamp 1669390400
transform 1 0 19824 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_169
timestamp 1669390400
transform 1 0 20272 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1669390400
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1669390400
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1669390400
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_456
timestamp 1669390400
transform 1 0 52416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_527
timestamp 1669390400
transform 1 0 60368 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1669390400
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_598
timestamp 1669390400
transform 1 0 68320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1669390400
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_605
timestamp 1669390400
transform 1 0 69104 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_669
timestamp 1669390400
transform 1 0 76272 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1669390400
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_676
timestamp 1669390400
transform 1 0 77056 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_684
timestamp 1669390400
transform 1 0 77952 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_20
timestamp 1669390400
transform 1 0 3584 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_24
timestamp 1669390400
transform 1 0 4032 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_28
timestamp 1669390400
transform 1 0 4480 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_32
timestamp 1669390400
transform 1 0 4928 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_36
timestamp 1669390400
transform 1 0 5376 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_42
timestamp 1669390400
transform 1 0 6048 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_46
timestamp 1669390400
transform 1 0 6496 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_50
timestamp 1669390400
transform 1 0 6944 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_54
timestamp 1669390400
transform 1 0 7392 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_58
timestamp 1669390400
transform 1 0 7840 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_62
timestamp 1669390400
transform 1 0 8288 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_66
timestamp 1669390400
transform 1 0 8736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1669390400
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_76
timestamp 1669390400
transform 1 0 9856 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_82
timestamp 1669390400
transform 1 0 10528 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_86
timestamp 1669390400
transform 1 0 10976 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_90
timestamp 1669390400
transform 1 0 11424 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_94
timestamp 1669390400
transform 1 0 11872 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_100
timestamp 1669390400
transform 1 0 12544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_106
timestamp 1669390400
transform 1 0 13216 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_110
timestamp 1669390400
transform 1 0 13664 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_112
timestamp 1669390400
transform 1 0 13888 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_115
timestamp 1669390400
transform 1 0 14224 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_119
timestamp 1669390400
transform 1 0 14672 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_122
timestamp 1669390400
transform 1 0 15008 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_124
timestamp 1669390400
transform 1 0 15232 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_127
timestamp 1669390400
transform 1 0 15568 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_131
timestamp 1669390400
transform 1 0 16016 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_133
timestamp 1669390400
transform 1 0 16240 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_136
timestamp 1669390400
transform 1 0 16576 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_140
timestamp 1669390400
transform 1 0 17024 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_147
timestamp 1669390400
transform 1 0 17808 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_151
timestamp 1669390400
transform 1 0 18256 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_155
timestamp 1669390400
transform 1 0 18704 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_159
timestamp 1669390400
transform 1 0 19152 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_191
timestamp 1669390400
transform 1 0 22736 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_207
timestamp 1669390400
transform 1 0 24528 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_211
timestamp 1669390400
transform 1 0 24976 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1669390400
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1669390400
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1669390400
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_421
timestamp 1669390400
transform 1 0 48496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1669390400
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1669390400
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1669390400
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_563
timestamp 1669390400
transform 1 0 64400 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_567
timestamp 1669390400
transform 1 0 64848 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1669390400
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_634
timestamp 1669390400
transform 1 0 72352 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1669390400
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_641
timestamp 1669390400
transform 1 0 73136 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_673
timestamp 1669390400
transform 1 0 76720 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_681
timestamp 1669390400
transform 1 0 77616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_685
timestamp 1669390400
transform 1 0 78064 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_687
timestamp 1669390400
transform 1 0 78288 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_8
timestamp 1669390400
transform 1 0 2240 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_12
timestamp 1669390400
transform 1 0 2688 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_16
timestamp 1669390400
transform 1 0 3136 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_20
timestamp 1669390400
transform 1 0 3584 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_24
timestamp 1669390400
transform 1 0 4032 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_28
timestamp 1669390400
transform 1 0 4480 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_32
timestamp 1669390400
transform 1 0 4928 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1669390400
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_41
timestamp 1669390400
transform 1 0 5936 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_45
timestamp 1669390400
transform 1 0 6384 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_49
timestamp 1669390400
transform 1 0 6832 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_53
timestamp 1669390400
transform 1 0 7280 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_55
timestamp 1669390400
transform 1 0 7504 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_58
timestamp 1669390400
transform 1 0 7840 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_62
timestamp 1669390400
transform 1 0 8288 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_66
timestamp 1669390400
transform 1 0 8736 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_70
timestamp 1669390400
transform 1 0 9184 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_74
timestamp 1669390400
transform 1 0 9632 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_76
timestamp 1669390400
transform 1 0 9856 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_79
timestamp 1669390400
transform 1 0 10192 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_85
timestamp 1669390400
transform 1 0 10864 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_89
timestamp 1669390400
transform 1 0 11312 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1669390400
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_108
timestamp 1669390400
transform 1 0 13440 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_111
timestamp 1669390400
transform 1 0 13776 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_113
timestamp 1669390400
transform 1 0 14000 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_116
timestamp 1669390400
transform 1 0 14336 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_120
timestamp 1669390400
transform 1 0 14784 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_126
timestamp 1669390400
transform 1 0 15456 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_130
timestamp 1669390400
transform 1 0 15904 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_132
timestamp 1669390400
transform 1 0 16128 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_135
timestamp 1669390400
transform 1 0 16464 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_139
timestamp 1669390400
transform 1 0 16912 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_143
timestamp 1669390400
transform 1 0 17360 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_147
timestamp 1669390400
transform 1 0 17808 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_149
timestamp 1669390400
transform 1 0 18032 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_152
timestamp 1669390400
transform 1 0 18368 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_156
timestamp 1669390400
transform 1 0 18816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_159
timestamp 1669390400
transform 1 0 19152 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_163
timestamp 1669390400
transform 1 0 19600 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_167
timestamp 1669390400
transform 1 0 20048 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_171
timestamp 1669390400
transform 1 0 20496 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_173
timestamp 1669390400
transform 1 0 20720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1669390400
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_179
timestamp 1669390400
transform 1 0 21392 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_185
timestamp 1669390400
transform 1 0 22064 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_193
timestamp 1669390400
transform 1 0 22960 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_197
timestamp 1669390400
transform 1 0 23408 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_201
timestamp 1669390400
transform 1 0 23856 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_233
timestamp 1669390400
transform 1 0 27440 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_241
timestamp 1669390400
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_245
timestamp 1669390400
transform 1 0 28784 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1669390400
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1669390400
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1669390400
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1669390400
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1669390400
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1669390400
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_456
timestamp 1669390400
transform 1 0 52416 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1669390400
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_463
timestamp 1669390400
transform 1 0 53200 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_527
timestamp 1669390400
transform 1 0 60368 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1669390400
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_598
timestamp 1669390400
transform 1 0 68320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1669390400
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_605
timestamp 1669390400
transform 1 0 69104 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_669
timestamp 1669390400
transform 1 0 76272 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_673
timestamp 1669390400
transform 1 0 76720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_676
timestamp 1669390400
transform 1 0 77056 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_684
timestamp 1669390400
transform 1 0 77952 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_6
timestamp 1669390400
transform 1 0 2016 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_10
timestamp 1669390400
transform 1 0 2464 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_14
timestamp 1669390400
transform 1 0 2912 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_18
timestamp 1669390400
transform 1 0 3360 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_22
timestamp 1669390400
transform 1 0 3808 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_26
timestamp 1669390400
transform 1 0 4256 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_30
timestamp 1669390400
transform 1 0 4704 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_34
timestamp 1669390400
transform 1 0 5152 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_38
timestamp 1669390400
transform 1 0 5600 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_42
timestamp 1669390400
transform 1 0 6048 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_46
timestamp 1669390400
transform 1 0 6496 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_50
timestamp 1669390400
transform 1 0 6944 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_54
timestamp 1669390400
transform 1 0 7392 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_58
timestamp 1669390400
transform 1 0 7840 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_62
timestamp 1669390400
transform 1 0 8288 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_66
timestamp 1669390400
transform 1 0 8736 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1669390400
transform 1 0 9184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_73
timestamp 1669390400
transform 1 0 9520 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_75
timestamp 1669390400
transform 1 0 9744 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_82
timestamp 1669390400
transform 1 0 10528 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_86
timestamp 1669390400
transform 1 0 10976 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_92
timestamp 1669390400
transform 1 0 11648 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_96
timestamp 1669390400
transform 1 0 12096 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_100
timestamp 1669390400
transform 1 0 12544 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_104
timestamp 1669390400
transform 1 0 12992 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_111
timestamp 1669390400
transform 1 0 13776 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_115
timestamp 1669390400
transform 1 0 14224 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_119
timestamp 1669390400
transform 1 0 14672 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_123
timestamp 1669390400
transform 1 0 15120 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_127
timestamp 1669390400
transform 1 0 15568 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_131
timestamp 1669390400
transform 1 0 16016 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_135
timestamp 1669390400
transform 1 0 16464 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1669390400
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_144
timestamp 1669390400
transform 1 0 17472 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_147
timestamp 1669390400
transform 1 0 17808 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_153
timestamp 1669390400
transform 1 0 18480 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_157
timestamp 1669390400
transform 1 0 18928 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_161
timestamp 1669390400
transform 1 0 19376 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_165
timestamp 1669390400
transform 1 0 19824 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_169
timestamp 1669390400
transform 1 0 20272 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_173
timestamp 1669390400
transform 1 0 20720 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_177
timestamp 1669390400
transform 1 0 21168 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_180
timestamp 1669390400
transform 1 0 21504 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_184
timestamp 1669390400
transform 1 0 21952 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_188
timestamp 1669390400
transform 1 0 22400 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_192
timestamp 1669390400
transform 1 0 22848 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_196
timestamp 1669390400
transform 1 0 23296 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_200
timestamp 1669390400
transform 1 0 23744 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_202
timestamp 1669390400
transform 1 0 23968 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_205
timestamp 1669390400
transform 1 0 24304 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_215
timestamp 1669390400
transform 1 0 25424 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_247
timestamp 1669390400
transform 1 0 29008 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_251
timestamp 1669390400
transform 1 0 29456 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_255
timestamp 1669390400
transform 1 0 29904 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_262
timestamp 1669390400
transform 1 0 30688 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_266
timestamp 1669390400
transform 1 0 31136 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_282
timestamp 1669390400
transform 1 0 32928 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1669390400
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1669390400
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_421
timestamp 1669390400
transform 1 0 48496 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1669390400
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1669390400
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_492
timestamp 1669390400
transform 1 0 56448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1669390400
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_499
timestamp 1669390400
transform 1 0 57232 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_563
timestamp 1669390400
transform 1 0 64400 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1669390400
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_570
timestamp 1669390400
transform 1 0 65184 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_634
timestamp 1669390400
transform 1 0 72352 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_638
timestamp 1669390400
transform 1 0 72800 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_641
timestamp 1669390400
transform 1 0 73136 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_673
timestamp 1669390400
transform 1 0 76720 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_681
timestamp 1669390400
transform 1 0 77616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_685
timestamp 1669390400
transform 1 0 78064 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_687
timestamp 1669390400
transform 1 0 78288 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_6
timestamp 1669390400
transform 1 0 2016 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_10
timestamp 1669390400
transform 1 0 2464 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_14
timestamp 1669390400
transform 1 0 2912 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_18
timestamp 1669390400
transform 1 0 3360 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_22
timestamp 1669390400
transform 1 0 3808 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_26
timestamp 1669390400
transform 1 0 4256 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_30
timestamp 1669390400
transform 1 0 4704 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_34
timestamp 1669390400
transform 1 0 5152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_37
timestamp 1669390400
transform 1 0 5488 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_39
timestamp 1669390400
transform 1 0 5712 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_42
timestamp 1669390400
transform 1 0 6048 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_46
timestamp 1669390400
transform 1 0 6496 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_50
timestamp 1669390400
transform 1 0 6944 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_54
timestamp 1669390400
transform 1 0 7392 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_56
timestamp 1669390400
transform 1 0 7616 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_59
timestamp 1669390400
transform 1 0 7952 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_65
timestamp 1669390400
transform 1 0 8624 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_69
timestamp 1669390400
transform 1 0 9072 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_73
timestamp 1669390400
transform 1 0 9520 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_77
timestamp 1669390400
transform 1 0 9968 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_81
timestamp 1669390400
transform 1 0 10416 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_89
timestamp 1669390400
transform 1 0 11312 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_93
timestamp 1669390400
transform 1 0 11760 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_97
timestamp 1669390400
transform 1 0 12208 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1669390400
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_108
timestamp 1669390400
transform 1 0 13440 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_117
timestamp 1669390400
transform 1 0 14448 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_121
timestamp 1669390400
transform 1 0 14896 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_125
timestamp 1669390400
transform 1 0 15344 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_135
timestamp 1669390400
transform 1 0 16464 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_139
timestamp 1669390400
transform 1 0 16912 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_143
timestamp 1669390400
transform 1 0 17360 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_147
timestamp 1669390400
transform 1 0 17808 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_151
timestamp 1669390400
transform 1 0 18256 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_157
timestamp 1669390400
transform 1 0 18928 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_161
timestamp 1669390400
transform 1 0 19376 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_165
timestamp 1669390400
transform 1 0 19824 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_171
timestamp 1669390400
transform 1 0 20496 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_175
timestamp 1669390400
transform 1 0 20944 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_179
timestamp 1669390400
transform 1 0 21392 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_181
timestamp 1669390400
transform 1 0 21616 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_184
timestamp 1669390400
transform 1 0 21952 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_188
timestamp 1669390400
transform 1 0 22400 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_192
timestamp 1669390400
transform 1 0 22848 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_196
timestamp 1669390400
transform 1 0 23296 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_200
timestamp 1669390400
transform 1 0 23744 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_202
timestamp 1669390400
transform 1 0 23968 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_205
timestamp 1669390400
transform 1 0 24304 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_209
timestamp 1669390400
transform 1 0 24752 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_212
timestamp 1669390400
transform 1 0 25088 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_216
timestamp 1669390400
transform 1 0 25536 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_220
timestamp 1669390400
transform 1 0 25984 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_236
timestamp 1669390400
transform 1 0 27776 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_244
timestamp 1669390400
transform 1 0 28672 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1669390400
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1669390400
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1669390400
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1669390400
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1669390400
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1669390400
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1669390400
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_456
timestamp 1669390400
transform 1 0 52416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1669390400
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_463
timestamp 1669390400
transform 1 0 53200 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_527
timestamp 1669390400
transform 1 0 60368 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1669390400
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_598
timestamp 1669390400
transform 1 0 68320 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1669390400
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_605
timestamp 1669390400
transform 1 0 69104 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_669
timestamp 1669390400
transform 1 0 76272 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1669390400
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_676
timestamp 1669390400
transform 1 0 77056 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_684
timestamp 1669390400
transform 1 0 77952 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_6
timestamp 1669390400
transform 1 0 2016 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_10
timestamp 1669390400
transform 1 0 2464 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_14
timestamp 1669390400
transform 1 0 2912 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_18
timestamp 1669390400
transform 1 0 3360 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_22
timestamp 1669390400
transform 1 0 3808 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_26
timestamp 1669390400
transform 1 0 4256 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_30
timestamp 1669390400
transform 1 0 4704 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_34
timestamp 1669390400
transform 1 0 5152 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_38
timestamp 1669390400
transform 1 0 5600 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_42
timestamp 1669390400
transform 1 0 6048 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_46
timestamp 1669390400
transform 1 0 6496 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_50
timestamp 1669390400
transform 1 0 6944 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_54
timestamp 1669390400
transform 1 0 7392 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_58
timestamp 1669390400
transform 1 0 7840 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_62
timestamp 1669390400
transform 1 0 8288 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_66
timestamp 1669390400
transform 1 0 8736 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_70
timestamp 1669390400
transform 1 0 9184 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_73
timestamp 1669390400
transform 1 0 9520 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_79
timestamp 1669390400
transform 1 0 10192 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_89
timestamp 1669390400
transform 1 0 11312 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_99
timestamp 1669390400
transform 1 0 12432 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_103
timestamp 1669390400
transform 1 0 12880 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_114
timestamp 1669390400
transform 1 0 14112 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_118
timestamp 1669390400
transform 1 0 14560 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_125
timestamp 1669390400
transform 1 0 15344 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_133
timestamp 1669390400
transform 1 0 16240 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_140
timestamp 1669390400
transform 1 0 17024 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_144
timestamp 1669390400
transform 1 0 17472 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_146
timestamp 1669390400
transform 1 0 17696 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_155
timestamp 1669390400
transform 1 0 18704 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_159
timestamp 1669390400
transform 1 0 19152 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_162
timestamp 1669390400
transform 1 0 19488 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_166
timestamp 1669390400
transform 1 0 19936 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_170
timestamp 1669390400
transform 1 0 20384 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_174
timestamp 1669390400
transform 1 0 20832 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_178
timestamp 1669390400
transform 1 0 21280 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_182
timestamp 1669390400
transform 1 0 21728 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_188
timestamp 1669390400
transform 1 0 22400 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_190
timestamp 1669390400
transform 1 0 22624 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_193
timestamp 1669390400
transform 1 0 22960 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_197
timestamp 1669390400
transform 1 0 23408 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_201
timestamp 1669390400
transform 1 0 23856 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_203
timestamp 1669390400
transform 1 0 24080 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_206
timestamp 1669390400
transform 1 0 24416 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_210
timestamp 1669390400
transform 1 0 24864 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1669390400
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_215
timestamp 1669390400
transform 1 0 25424 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_218
timestamp 1669390400
transform 1 0 25760 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_220
timestamp 1669390400
transform 1 0 25984 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_223
timestamp 1669390400
transform 1 0 26320 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_227
timestamp 1669390400
transform 1 0 26768 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_231
timestamp 1669390400
transform 1 0 27216 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_233
timestamp 1669390400
transform 1 0 27440 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_236
timestamp 1669390400
transform 1 0 27776 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_243
timestamp 1669390400
transform 1 0 28560 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_247
timestamp 1669390400
transform 1 0 29008 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1669390400
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1669390400
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1669390400
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1669390400
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1669390400
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1669390400
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1669390400
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_492
timestamp 1669390400
transform 1 0 56448 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1669390400
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_499
timestamp 1669390400
transform 1 0 57232 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_563
timestamp 1669390400
transform 1 0 64400 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1669390400
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_570
timestamp 1669390400
transform 1 0 65184 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_634
timestamp 1669390400
transform 1 0 72352 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1669390400
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_641
timestamp 1669390400
transform 1 0 73136 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_673
timestamp 1669390400
transform 1 0 76720 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_681
timestamp 1669390400
transform 1 0 77616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_685
timestamp 1669390400
transform 1 0 78064 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_687
timestamp 1669390400
transform 1 0 78288 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_6
timestamp 1669390400
transform 1 0 2016 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_10
timestamp 1669390400
transform 1 0 2464 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_14
timestamp 1669390400
transform 1 0 2912 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_18
timestamp 1669390400
transform 1 0 3360 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_22
timestamp 1669390400
transform 1 0 3808 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_26
timestamp 1669390400
transform 1 0 4256 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_30
timestamp 1669390400
transform 1 0 4704 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_34
timestamp 1669390400
transform 1 0 5152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_37
timestamp 1669390400
transform 1 0 5488 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_43
timestamp 1669390400
transform 1 0 6160 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_47
timestamp 1669390400
transform 1 0 6608 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_51
timestamp 1669390400
transform 1 0 7056 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_55
timestamp 1669390400
transform 1 0 7504 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_59
timestamp 1669390400
transform 1 0 7952 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_63
timestamp 1669390400
transform 1 0 8400 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_67
timestamp 1669390400
transform 1 0 8848 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_74
timestamp 1669390400
transform 1 0 9632 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_84
timestamp 1669390400
transform 1 0 10752 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_99
timestamp 1669390400
transform 1 0 12432 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1669390400
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_108
timestamp 1669390400
transform 1 0 13440 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_121
timestamp 1669390400
transform 1 0 14896 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_123
timestamp 1669390400
transform 1 0 15120 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_126
timestamp 1669390400
transform 1 0 15456 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_141
timestamp 1669390400
transform 1 0 17136 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_160
timestamp 1669390400
transform 1 0 19264 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_167
timestamp 1669390400
transform 1 0 20048 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_169
timestamp 1669390400
transform 1 0 20272 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_172
timestamp 1669390400
transform 1 0 20608 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1669390400
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_179
timestamp 1669390400
transform 1 0 21392 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_189
timestamp 1669390400
transform 1 0 22512 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_195
timestamp 1669390400
transform 1 0 23184 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_201
timestamp 1669390400
transform 1 0 23856 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_208
timestamp 1669390400
transform 1 0 24640 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_215
timestamp 1669390400
transform 1 0 25424 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_221
timestamp 1669390400
transform 1 0 26096 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_225
timestamp 1669390400
transform 1 0 26544 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_229
timestamp 1669390400
transform 1 0 26992 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_233
timestamp 1669390400
transform 1 0 27440 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_237
timestamp 1669390400
transform 1 0 27888 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_243
timestamp 1669390400
transform 1 0 28560 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1669390400
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_250
timestamp 1669390400
transform 1 0 29344 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_257
timestamp 1669390400
transform 1 0 30128 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_289
timestamp 1669390400
transform 1 0 33712 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_305
timestamp 1669390400
transform 1 0 35504 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_313
timestamp 1669390400
transform 1 0 36400 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_317
timestamp 1669390400
transform 1 0 36848 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1669390400
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1669390400
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1669390400
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1669390400
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_456
timestamp 1669390400
transform 1 0 52416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1669390400
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_463
timestamp 1669390400
transform 1 0 53200 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_527
timestamp 1669390400
transform 1 0 60368 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_531
timestamp 1669390400
transform 1 0 60816 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_598
timestamp 1669390400
transform 1 0 68320 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1669390400
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_605
timestamp 1669390400
transform 1 0 69104 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_669
timestamp 1669390400
transform 1 0 76272 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1669390400
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_676
timestamp 1669390400
transform 1 0 77056 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_684
timestamp 1669390400
transform 1 0 77952 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_6
timestamp 1669390400
transform 1 0 2016 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_10
timestamp 1669390400
transform 1 0 2464 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_14
timestamp 1669390400
transform 1 0 2912 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_18
timestamp 1669390400
transform 1 0 3360 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_22
timestamp 1669390400
transform 1 0 3808 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_26
timestamp 1669390400
transform 1 0 4256 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_30
timestamp 1669390400
transform 1 0 4704 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_34
timestamp 1669390400
transform 1 0 5152 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_38
timestamp 1669390400
transform 1 0 5600 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_42
timestamp 1669390400
transform 1 0 6048 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_46
timestamp 1669390400
transform 1 0 6496 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_50
timestamp 1669390400
transform 1 0 6944 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_54
timestamp 1669390400
transform 1 0 7392 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_58
timestamp 1669390400
transform 1 0 7840 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_68
timestamp 1669390400
transform 1 0 8960 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1669390400
transform 1 0 9184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_73
timestamp 1669390400
transform 1 0 9520 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_88
timestamp 1669390400
transform 1 0 11200 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_92
timestamp 1669390400
transform 1 0 11648 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_102
timestamp 1669390400
transform 1 0 12768 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_117
timestamp 1669390400
transform 1 0 14448 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_119
timestamp 1669390400
transform 1 0 14672 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_130
timestamp 1669390400
transform 1 0 15904 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_132
timestamp 1669390400
transform 1 0 16128 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1669390400
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_144
timestamp 1669390400
transform 1 0 17472 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_155
timestamp 1669390400
transform 1 0 18704 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_165
timestamp 1669390400
transform 1 0 19824 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_172
timestamp 1669390400
transform 1 0 20608 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_188
timestamp 1669390400
transform 1 0 22400 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_198
timestamp 1669390400
transform 1 0 23520 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_206
timestamp 1669390400
transform 1 0 24416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1669390400
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_215
timestamp 1669390400
transform 1 0 25424 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_221
timestamp 1669390400
transform 1 0 26096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_233
timestamp 1669390400
transform 1 0 27440 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_237
timestamp 1669390400
transform 1 0 27888 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_241
timestamp 1669390400
transform 1 0 28336 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_244
timestamp 1669390400
transform 1 0 28672 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_248
timestamp 1669390400
transform 1 0 29120 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_280
timestamp 1669390400
transform 1 0 32704 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1669390400
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1669390400
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1669390400
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1669390400
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1669390400
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_492
timestamp 1669390400
transform 1 0 56448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1669390400
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_499
timestamp 1669390400
transform 1 0 57232 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_563
timestamp 1669390400
transform 1 0 64400 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1669390400
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_570
timestamp 1669390400
transform 1 0 65184 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_634
timestamp 1669390400
transform 1 0 72352 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1669390400
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_641
timestamp 1669390400
transform 1 0 73136 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_673
timestamp 1669390400
transform 1 0 76720 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_681
timestamp 1669390400
transform 1 0 77616 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_685
timestamp 1669390400
transform 1 0 78064 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_687
timestamp 1669390400
transform 1 0 78288 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_6
timestamp 1669390400
transform 1 0 2016 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_10
timestamp 1669390400
transform 1 0 2464 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_14
timestamp 1669390400
transform 1 0 2912 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_18
timestamp 1669390400
transform 1 0 3360 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_22
timestamp 1669390400
transform 1 0 3808 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_26
timestamp 1669390400
transform 1 0 4256 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_30
timestamp 1669390400
transform 1 0 4704 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_34
timestamp 1669390400
transform 1 0 5152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_37
timestamp 1669390400
transform 1 0 5488 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_39
timestamp 1669390400
transform 1 0 5712 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_63
timestamp 1669390400
transform 1 0 8400 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_69
timestamp 1669390400
transform 1 0 9072 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_81
timestamp 1669390400
transform 1 0 10416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_87
timestamp 1669390400
transform 1 0 11088 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_104
timestamp 1669390400
transform 1 0 12992 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_108
timestamp 1669390400
transform 1 0 13440 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_122
timestamp 1669390400
transform 1 0 15008 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_134
timestamp 1669390400
transform 1 0 16352 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_148
timestamp 1669390400
transform 1 0 17920 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_158
timestamp 1669390400
transform 1 0 19040 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_160
timestamp 1669390400
transform 1 0 19264 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_175
timestamp 1669390400
transform 1 0 20944 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_179
timestamp 1669390400
transform 1 0 21392 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_191
timestamp 1669390400
transform 1 0 22736 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_193
timestamp 1669390400
transform 1 0 22960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_196
timestamp 1669390400
transform 1 0 23296 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_207
timestamp 1669390400
transform 1 0 24528 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_221
timestamp 1669390400
transform 1 0 26096 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_230
timestamp 1669390400
transform 1 0 27104 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_244
timestamp 1669390400
transform 1 0 28672 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_250
timestamp 1669390400
transform 1 0 29344 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_256
timestamp 1669390400
transform 1 0 30016 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_260
timestamp 1669390400
transform 1 0 30464 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_292
timestamp 1669390400
transform 1 0 34048 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_308
timestamp 1669390400
transform 1 0 35840 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_316
timestamp 1669390400
transform 1 0 36736 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1669390400
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1669390400
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1669390400
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1669390400
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1669390400
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_456
timestamp 1669390400
transform 1 0 52416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1669390400
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1669390400
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_527
timestamp 1669390400
transform 1 0 60368 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1669390400
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_598
timestamp 1669390400
transform 1 0 68320 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1669390400
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_605
timestamp 1669390400
transform 1 0 69104 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_669
timestamp 1669390400
transform 1 0 76272 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1669390400
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_676
timestamp 1669390400
transform 1 0 77056 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_684
timestamp 1669390400
transform 1 0 77952 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_5
timestamp 1669390400
transform 1 0 1904 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_9
timestamp 1669390400
transform 1 0 2352 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_13
timestamp 1669390400
transform 1 0 2800 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_17
timestamp 1669390400
transform 1 0 3248 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_21
timestamp 1669390400
transform 1 0 3696 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_25
timestamp 1669390400
transform 1 0 4144 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_29
timestamp 1669390400
transform 1 0 4592 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_33
timestamp 1669390400
transform 1 0 5040 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_39
timestamp 1669390400
transform 1 0 5712 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_43
timestamp 1669390400
transform 1 0 6160 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_46
timestamp 1669390400
transform 1 0 6496 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_50
timestamp 1669390400
transform 1 0 6944 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_57
timestamp 1669390400
transform 1 0 7728 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_67
timestamp 1669390400
transform 1 0 8848 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_73
timestamp 1669390400
transform 1 0 9520 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_83
timestamp 1669390400
transform 1 0 10640 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_103
timestamp 1669390400
transform 1 0 12880 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_129
timestamp 1669390400
transform 1 0 15792 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_140
timestamp 1669390400
transform 1 0 17024 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_144
timestamp 1669390400
transform 1 0 17472 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_156
timestamp 1669390400
transform 1 0 18816 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_160
timestamp 1669390400
transform 1 0 19264 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_173
timestamp 1669390400
transform 1 0 20720 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_186
timestamp 1669390400
transform 1 0 22176 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_194
timestamp 1669390400
transform 1 0 23072 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_207
timestamp 1669390400
transform 1 0 24528 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_209
timestamp 1669390400
transform 1 0 24752 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1669390400
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_215
timestamp 1669390400
transform 1 0 25424 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_228
timestamp 1669390400
transform 1 0 26880 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_239
timestamp 1669390400
transform 1 0 28112 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_243
timestamp 1669390400
transform 1 0 28560 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_256
timestamp 1669390400
transform 1 0 30016 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_263
timestamp 1669390400
transform 1 0 30800 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_267
timestamp 1669390400
transform 1 0 31248 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1669390400
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1669390400
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1669390400
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1669390400
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1669390400
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1669390400
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_492
timestamp 1669390400
transform 1 0 56448 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1669390400
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_499
timestamp 1669390400
transform 1 0 57232 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_563
timestamp 1669390400
transform 1 0 64400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1669390400
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_570
timestamp 1669390400
transform 1 0 65184 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_634
timestamp 1669390400
transform 1 0 72352 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_638
timestamp 1669390400
transform 1 0 72800 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_641
timestamp 1669390400
transform 1 0 73136 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_673
timestamp 1669390400
transform 1 0 76720 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_681
timestamp 1669390400
transform 1 0 77616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_685
timestamp 1669390400
transform 1 0 78064 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_687
timestamp 1669390400
transform 1 0 78288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_8
timestamp 1669390400
transform 1 0 2240 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_12
timestamp 1669390400
transform 1 0 2688 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_20
timestamp 1669390400
transform 1 0 3584 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_26
timestamp 1669390400
transform 1 0 4256 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_30
timestamp 1669390400
transform 1 0 4704 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1669390400
transform 1 0 5152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_37
timestamp 1669390400
transform 1 0 5488 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_41
timestamp 1669390400
transform 1 0 5936 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_45
timestamp 1669390400
transform 1 0 6384 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_51
timestamp 1669390400
transform 1 0 7056 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_57
timestamp 1669390400
transform 1 0 7728 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_65
timestamp 1669390400
transform 1 0 8624 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_73
timestamp 1669390400
transform 1 0 9520 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_98
timestamp 1669390400
transform 1 0 12320 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1669390400
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_108
timestamp 1669390400
transform 1 0 13440 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_138
timestamp 1669390400
transform 1 0 16800 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_150
timestamp 1669390400
transform 1 0 18144 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_157
timestamp 1669390400
transform 1 0 18928 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_171
timestamp 1669390400
transform 1 0 20496 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_173
timestamp 1669390400
transform 1 0 20720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1669390400
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_179
timestamp 1669390400
transform 1 0 21392 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_181
timestamp 1669390400
transform 1 0 21616 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_194
timestamp 1669390400
transform 1 0 23072 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_225
timestamp 1669390400
transform 1 0 26544 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_235
timestamp 1669390400
transform 1 0 27664 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1669390400
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_250
timestamp 1669390400
transform 1 0 29344 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_257
timestamp 1669390400
transform 1 0 30128 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_259
timestamp 1669390400
transform 1 0 30352 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_272
timestamp 1669390400
transform 1 0 31808 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_276
timestamp 1669390400
transform 1 0 32256 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_308
timestamp 1669390400
transform 1 0 35840 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_316
timestamp 1669390400
transform 1 0 36736 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1669390400
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1669390400
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1669390400
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1669390400
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1669390400
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_456
timestamp 1669390400
transform 1 0 52416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1669390400
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1669390400
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_527
timestamp 1669390400
transform 1 0 60368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1669390400
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_598
timestamp 1669390400
transform 1 0 68320 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1669390400
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_605
timestamp 1669390400
transform 1 0 69104 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_669
timestamp 1669390400
transform 1 0 76272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1669390400
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_676
timestamp 1669390400
transform 1 0 77056 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_684
timestamp 1669390400
transform 1 0 77952 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_6
timestamp 1669390400
transform 1 0 2016 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_10
timestamp 1669390400
transform 1 0 2464 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_14
timestamp 1669390400
transform 1 0 2912 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_18
timestamp 1669390400
transform 1 0 3360 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_22
timestamp 1669390400
transform 1 0 3808 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_26
timestamp 1669390400
transform 1 0 4256 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_30
timestamp 1669390400
transform 1 0 4704 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_34
timestamp 1669390400
transform 1 0 5152 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_38
timestamp 1669390400
transform 1 0 5600 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_42
timestamp 1669390400
transform 1 0 6048 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_50
timestamp 1669390400
transform 1 0 6944 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_58
timestamp 1669390400
transform 1 0 7840 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1669390400
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_73
timestamp 1669390400
transform 1 0 9520 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_75
timestamp 1669390400
transform 1 0 9744 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_84
timestamp 1669390400
transform 1 0 10752 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_88
timestamp 1669390400
transform 1 0 11200 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_118
timestamp 1669390400
transform 1 0 14560 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_132
timestamp 1669390400
transform 1 0 16128 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_134
timestamp 1669390400
transform 1 0 16352 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1669390400
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_144
timestamp 1669390400
transform 1 0 17472 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_155
timestamp 1669390400
transform 1 0 18704 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_188
timestamp 1669390400
transform 1 0 22400 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_192
timestamp 1669390400
transform 1 0 22848 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_207
timestamp 1669390400
transform 1 0 24528 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_209
timestamp 1669390400
transform 1 0 24752 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1669390400
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_215
timestamp 1669390400
transform 1 0 25424 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_224
timestamp 1669390400
transform 1 0 26432 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_231
timestamp 1669390400
transform 1 0 27216 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_239
timestamp 1669390400
transform 1 0 28112 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_245
timestamp 1669390400
transform 1 0 28784 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_264
timestamp 1669390400
transform 1 0 30912 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_271
timestamp 1669390400
transform 1 0 31696 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_275
timestamp 1669390400
transform 1 0 32144 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_279
timestamp 1669390400
transform 1 0 32592 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1669390400
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1669390400
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1669390400
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_421
timestamp 1669390400
transform 1 0 48496 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1669390400
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1669390400
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_492
timestamp 1669390400
transform 1 0 56448 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1669390400
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_499
timestamp 1669390400
transform 1 0 57232 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_563
timestamp 1669390400
transform 1 0 64400 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1669390400
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_570
timestamp 1669390400
transform 1 0 65184 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_634
timestamp 1669390400
transform 1 0 72352 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1669390400
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_641
timestamp 1669390400
transform 1 0 73136 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_673
timestamp 1669390400
transform 1 0 76720 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_681
timestamp 1669390400
transform 1 0 77616 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_685
timestamp 1669390400
transform 1 0 78064 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_687
timestamp 1669390400
transform 1 0 78288 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_6
timestamp 1669390400
transform 1 0 2016 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_10
timestamp 1669390400
transform 1 0 2464 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_14
timestamp 1669390400
transform 1 0 2912 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_18
timestamp 1669390400
transform 1 0 3360 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_22
timestamp 1669390400
transform 1 0 3808 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_26
timestamp 1669390400
transform 1 0 4256 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_30
timestamp 1669390400
transform 1 0 4704 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1669390400
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_37
timestamp 1669390400
transform 1 0 5488 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_39
timestamp 1669390400
transform 1 0 5712 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_45
timestamp 1669390400
transform 1 0 6384 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_55
timestamp 1669390400
transform 1 0 7504 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_65
timestamp 1669390400
transform 1 0 8624 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_75
timestamp 1669390400
transform 1 0 9744 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_85
timestamp 1669390400
transform 1 0 10864 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_95
timestamp 1669390400
transform 1 0 11984 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1669390400
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_108
timestamp 1669390400
transform 1 0 13440 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_119
timestamp 1669390400
transform 1 0 14672 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_139
timestamp 1669390400
transform 1 0 16912 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_143
timestamp 1669390400
transform 1 0 17360 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1669390400
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_179
timestamp 1669390400
transform 1 0 21392 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_192
timestamp 1669390400
transform 1 0 22848 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_203
timestamp 1669390400
transform 1 0 24080 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_210
timestamp 1669390400
transform 1 0 24864 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_241
timestamp 1669390400
transform 1 0 28336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1669390400
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_250
timestamp 1669390400
transform 1 0 29344 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_257
timestamp 1669390400
transform 1 0 30128 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_264
timestamp 1669390400
transform 1 0 30912 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_268
timestamp 1669390400
transform 1 0 31360 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_274
timestamp 1669390400
transform 1 0 32032 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_281
timestamp 1669390400
transform 1 0 32816 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_285
timestamp 1669390400
transform 1 0 33264 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_289
timestamp 1669390400
transform 1 0 33712 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_293
timestamp 1669390400
transform 1 0 34160 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_297
timestamp 1669390400
transform 1 0 34608 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_313
timestamp 1669390400
transform 1 0 36400 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_317
timestamp 1669390400
transform 1 0 36848 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1669390400
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1669390400
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1669390400
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1669390400
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_456
timestamp 1669390400
transform 1 0 52416 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1669390400
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_463
timestamp 1669390400
transform 1 0 53200 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_527
timestamp 1669390400
transform 1 0 60368 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1669390400
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_598
timestamp 1669390400
transform 1 0 68320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1669390400
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_605
timestamp 1669390400
transform 1 0 69104 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_669
timestamp 1669390400
transform 1 0 76272 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_673
timestamp 1669390400
transform 1 0 76720 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_676
timestamp 1669390400
transform 1 0 77056 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_684
timestamp 1669390400
transform 1 0 77952 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_4
timestamp 1669390400
transform 1 0 1792 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_7
timestamp 1669390400
transform 1 0 2128 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_11
timestamp 1669390400
transform 1 0 2576 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_15
timestamp 1669390400
transform 1 0 3024 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_19
timestamp 1669390400
transform 1 0 3472 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_23
timestamp 1669390400
transform 1 0 3920 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_29
timestamp 1669390400
transform 1 0 4592 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_37
timestamp 1669390400
transform 1 0 5488 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_70
timestamp 1669390400
transform 1 0 9184 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_73
timestamp 1669390400
transform 1 0 9520 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_78
timestamp 1669390400
transform 1 0 10080 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_88
timestamp 1669390400
transform 1 0 11200 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_140
timestamp 1669390400
transform 1 0 17024 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_144
timestamp 1669390400
transform 1 0 17472 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_156
timestamp 1669390400
transform 1 0 18816 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_208
timestamp 1669390400
transform 1 0 24640 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1669390400
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_215
timestamp 1669390400
transform 1 0 25424 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_225
timestamp 1669390400
transform 1 0 26544 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_235
timestamp 1669390400
transform 1 0 27664 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_239
timestamp 1669390400
transform 1 0 28112 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_259
timestamp 1669390400
transform 1 0 30352 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_274
timestamp 1669390400
transform 1 0 32032 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1669390400
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_286
timestamp 1669390400
transform 1 0 33376 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_289
timestamp 1669390400
transform 1 0 33712 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_293
timestamp 1669390400
transform 1 0 34160 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_297
timestamp 1669390400
transform 1 0 34608 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_301
timestamp 1669390400
transform 1 0 35056 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_305
timestamp 1669390400
transform 1 0 35504 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_337
timestamp 1669390400
transform 1 0 39088 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_353
timestamp 1669390400
transform 1 0 40880 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1669390400
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1669390400
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1669390400
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_492
timestamp 1669390400
transform 1 0 56448 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1669390400
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1669390400
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_563
timestamp 1669390400
transform 1 0 64400 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1669390400
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_570
timestamp 1669390400
transform 1 0 65184 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_634
timestamp 1669390400
transform 1 0 72352 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1669390400
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_641
timestamp 1669390400
transform 1 0 73136 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_673
timestamp 1669390400
transform 1 0 76720 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_681
timestamp 1669390400
transform 1 0 77616 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_685
timestamp 1669390400
transform 1 0 78064 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_687
timestamp 1669390400
transform 1 0 78288 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_6
timestamp 1669390400
transform 1 0 2016 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_10
timestamp 1669390400
transform 1 0 2464 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_14
timestamp 1669390400
transform 1 0 2912 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_18
timestamp 1669390400
transform 1 0 3360 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_22
timestamp 1669390400
transform 1 0 3808 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_26
timestamp 1669390400
transform 1 0 4256 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_30
timestamp 1669390400
transform 1 0 4704 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_34
timestamp 1669390400
transform 1 0 5152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_37
timestamp 1669390400
transform 1 0 5488 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_47
timestamp 1669390400
transform 1 0 6608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_53
timestamp 1669390400
transform 1 0 7280 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_63
timestamp 1669390400
transform 1 0 8400 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_88
timestamp 1669390400
transform 1 0 11200 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_95
timestamp 1669390400
transform 1 0 11984 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1669390400
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_108
timestamp 1669390400
transform 1 0 13440 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_138
timestamp 1669390400
transform 1 0 16800 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_169
timestamp 1669390400
transform 1 0 20272 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1669390400
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_179
timestamp 1669390400
transform 1 0 21392 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_183
timestamp 1669390400
transform 1 0 21840 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_214
timestamp 1669390400
transform 1 0 25312 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_224
timestamp 1669390400
transform 1 0 26432 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_234
timestamp 1669390400
transform 1 0 27552 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_236
timestamp 1669390400
transform 1 0 27776 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1669390400
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_250
timestamp 1669390400
transform 1 0 29344 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_259
timestamp 1669390400
transform 1 0 30352 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_265
timestamp 1669390400
transform 1 0 31024 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_269
timestamp 1669390400
transform 1 0 31472 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_276
timestamp 1669390400
transform 1 0 32256 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_283
timestamp 1669390400
transform 1 0 33040 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_289
timestamp 1669390400
transform 1 0 33712 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_293
timestamp 1669390400
transform 1 0 34160 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_297
timestamp 1669390400
transform 1 0 34608 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_301
timestamp 1669390400
transform 1 0 35056 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_305
timestamp 1669390400
transform 1 0 35504 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_309
timestamp 1669390400
transform 1 0 35952 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_313
timestamp 1669390400
transform 1 0 36400 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_317
timestamp 1669390400
transform 1 0 36848 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1669390400
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1669390400
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1669390400
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1669390400
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1669390400
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1669390400
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1669390400
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_527
timestamp 1669390400
transform 1 0 60368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1669390400
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1669390400
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1669390400
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1669390400
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_605
timestamp 1669390400
transform 1 0 69104 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_669
timestamp 1669390400
transform 1 0 76272 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1669390400
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_676
timestamp 1669390400
transform 1 0 77056 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_684
timestamp 1669390400
transform 1 0 77952 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_12
timestamp 1669390400
transform 1 0 2688 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_16
timestamp 1669390400
transform 1 0 3136 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_20
timestamp 1669390400
transform 1 0 3584 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_24
timestamp 1669390400
transform 1 0 4032 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_28
timestamp 1669390400
transform 1 0 4480 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_32
timestamp 1669390400
transform 1 0 4928 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_42
timestamp 1669390400
transform 1 0 6048 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_46
timestamp 1669390400
transform 1 0 6496 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_49
timestamp 1669390400
transform 1 0 6832 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_57
timestamp 1669390400
transform 1 0 7728 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_68
timestamp 1669390400
transform 1 0 8960 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_70
timestamp 1669390400
transform 1 0 9184 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_73
timestamp 1669390400
transform 1 0 9520 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_75
timestamp 1669390400
transform 1 0 9744 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_105
timestamp 1669390400
transform 1 0 13104 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_138
timestamp 1669390400
transform 1 0 16800 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_144
timestamp 1669390400
transform 1 0 17472 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_159
timestamp 1669390400
transform 1 0 19152 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_161
timestamp 1669390400
transform 1 0 19376 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_164
timestamp 1669390400
transform 1 0 19712 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_197
timestamp 1669390400
transform 1 0 23408 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_207
timestamp 1669390400
transform 1 0 24528 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_209
timestamp 1669390400
transform 1 0 24752 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1669390400
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_215
timestamp 1669390400
transform 1 0 25424 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_245
timestamp 1669390400
transform 1 0 28784 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_256
timestamp 1669390400
transform 1 0 30016 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_258
timestamp 1669390400
transform 1 0 30240 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_271
timestamp 1669390400
transform 1 0 31696 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_281
timestamp 1669390400
transform 1 0 32816 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1669390400
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_286
timestamp 1669390400
transform 1 0 33376 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_295
timestamp 1669390400
transform 1 0 34384 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_299
timestamp 1669390400
transform 1 0 34832 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_303
timestamp 1669390400
transform 1 0 35280 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_307
timestamp 1669390400
transform 1 0 35728 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_311
timestamp 1669390400
transform 1 0 36176 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_315
timestamp 1669390400
transform 1 0 36624 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_319
timestamp 1669390400
transform 1 0 37072 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_323
timestamp 1669390400
transform 1 0 37520 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1669390400
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1669390400
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1669390400
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1669390400
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1669390400
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1669390400
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1669390400
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1669390400
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_570
timestamp 1669390400
transform 1 0 65184 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_634
timestamp 1669390400
transform 1 0 72352 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1669390400
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_641
timestamp 1669390400
transform 1 0 73136 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_673
timestamp 1669390400
transform 1 0 76720 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_681
timestamp 1669390400
transform 1 0 77616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_685
timestamp 1669390400
transform 1 0 78064 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_687
timestamp 1669390400
transform 1 0 78288 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_8
timestamp 1669390400
transform 1 0 2240 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_12
timestamp 1669390400
transform 1 0 2688 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_16
timestamp 1669390400
transform 1 0 3136 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_20
timestamp 1669390400
transform 1 0 3584 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_24
timestamp 1669390400
transform 1 0 4032 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1669390400
transform 1 0 5152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_37
timestamp 1669390400
transform 1 0 5488 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_49
timestamp 1669390400
transform 1 0 6832 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_56
timestamp 1669390400
transform 1 0 7616 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_89
timestamp 1669390400
transform 1 0 11312 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_95
timestamp 1669390400
transform 1 0 11984 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1669390400
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_108
timestamp 1669390400
transform 1 0 13440 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_121
timestamp 1669390400
transform 1 0 14896 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_173
timestamp 1669390400
transform 1 0 20720 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_179
timestamp 1669390400
transform 1 0 21392 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_209
timestamp 1669390400
transform 1 0 24752 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_226
timestamp 1669390400
transform 1 0 26656 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_240
timestamp 1669390400
transform 1 0 28224 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_246
timestamp 1669390400
transform 1 0 28896 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_250
timestamp 1669390400
transform 1 0 29344 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_261
timestamp 1669390400
transform 1 0 30576 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_263
timestamp 1669390400
transform 1 0 30800 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_276
timestamp 1669390400
transform 1 0 32256 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_284
timestamp 1669390400
transform 1 0 33152 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_291
timestamp 1669390400
transform 1 0 33936 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_295
timestamp 1669390400
transform 1 0 34384 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_299
timestamp 1669390400
transform 1 0 34832 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_303
timestamp 1669390400
transform 1 0 35280 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_307
timestamp 1669390400
transform 1 0 35728 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_311
timestamp 1669390400
transform 1 0 36176 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_315
timestamp 1669390400
transform 1 0 36624 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_321
timestamp 1669390400
transform 1 0 37296 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_324
timestamp 1669390400
transform 1 0 37632 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_328
timestamp 1669390400
transform 1 0 38080 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_332
timestamp 1669390400
transform 1 0 38528 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_364
timestamp 1669390400
transform 1 0 42112 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_380
timestamp 1669390400
transform 1 0 43904 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_388
timestamp 1669390400
transform 1 0 44800 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1669390400
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1669390400
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1669390400
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1669390400
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1669390400
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1669390400
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1669390400
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1669390400
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_605
timestamp 1669390400
transform 1 0 69104 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_669
timestamp 1669390400
transform 1 0 76272 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_673
timestamp 1669390400
transform 1 0 76720 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_676
timestamp 1669390400
transform 1 0 77056 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_684
timestamp 1669390400
transform 1 0 77952 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_6
timestamp 1669390400
transform 1 0 2016 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_10
timestamp 1669390400
transform 1 0 2464 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_14
timestamp 1669390400
transform 1 0 2912 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_28
timestamp 1669390400
transform 1 0 4480 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_30
timestamp 1669390400
transform 1 0 4704 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_33
timestamp 1669390400
transform 1 0 5040 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_43
timestamp 1669390400
transform 1 0 6160 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_68
timestamp 1669390400
transform 1 0 8960 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_70
timestamp 1669390400
transform 1 0 9184 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_73
timestamp 1669390400
transform 1 0 9520 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_76
timestamp 1669390400
transform 1 0 9856 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_88
timestamp 1669390400
transform 1 0 11200 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_140
timestamp 1669390400
transform 1 0 17024 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_144
timestamp 1669390400
transform 1 0 17472 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_156
timestamp 1669390400
transform 1 0 18816 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_208
timestamp 1669390400
transform 1 0 24640 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1669390400
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_215
timestamp 1669390400
transform 1 0 25424 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_224
timestamp 1669390400
transform 1 0 26432 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_238
timestamp 1669390400
transform 1 0 28000 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_272
timestamp 1669390400
transform 1 0 31808 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_274
timestamp 1669390400
transform 1 0 32032 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1669390400
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_286
timestamp 1669390400
transform 1 0 33376 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_295
timestamp 1669390400
transform 1 0 34384 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_299
timestamp 1669390400
transform 1 0 34832 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_303
timestamp 1669390400
transform 1 0 35280 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_307
timestamp 1669390400
transform 1 0 35728 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_311
timestamp 1669390400
transform 1 0 36176 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_315
timestamp 1669390400
transform 1 0 36624 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_319
timestamp 1669390400
transform 1 0 37072 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_323
timestamp 1669390400
transform 1 0 37520 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_327
timestamp 1669390400
transform 1 0 37968 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_331
timestamp 1669390400
transform 1 0 38416 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_347
timestamp 1669390400
transform 1 0 40208 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1669390400
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1669390400
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1669390400
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1669390400
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1669390400
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1669390400
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1669390400
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1669390400
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_570
timestamp 1669390400
transform 1 0 65184 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_634
timestamp 1669390400
transform 1 0 72352 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1669390400
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_641
timestamp 1669390400
transform 1 0 73136 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_673
timestamp 1669390400
transform 1 0 76720 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_681
timestamp 1669390400
transform 1 0 77616 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_685
timestamp 1669390400
transform 1 0 78064 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_687
timestamp 1669390400
transform 1 0 78288 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_4
timestamp 1669390400
transform 1 0 1792 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_7
timestamp 1669390400
transform 1 0 2128 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_11
timestamp 1669390400
transform 1 0 2576 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_15
timestamp 1669390400
transform 1 0 3024 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_19
timestamp 1669390400
transform 1 0 3472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_23
timestamp 1669390400
transform 1 0 3920 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_27
timestamp 1669390400
transform 1 0 4368 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1669390400
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_37
timestamp 1669390400
transform 1 0 5488 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_39
timestamp 1669390400
transform 1 0 5712 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_46
timestamp 1669390400
transform 1 0 6496 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_56
timestamp 1669390400
transform 1 0 7616 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_66
timestamp 1669390400
transform 1 0 8736 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_82
timestamp 1669390400
transform 1 0 10528 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_89
timestamp 1669390400
transform 1 0 11312 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_103
timestamp 1669390400
transform 1 0 12880 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1669390400
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_108
timestamp 1669390400
transform 1 0 13440 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_113
timestamp 1669390400
transform 1 0 14000 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_146
timestamp 1669390400
transform 1 0 17696 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_157
timestamp 1669390400
transform 1 0 18928 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_159
timestamp 1669390400
transform 1 0 19152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_166
timestamp 1669390400
transform 1 0 19936 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1669390400
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_179
timestamp 1669390400
transform 1 0 21392 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_209
timestamp 1669390400
transform 1 0 24752 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_211
timestamp 1669390400
transform 1 0 24976 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_214
timestamp 1669390400
transform 1 0 25312 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1669390400
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_250
timestamp 1669390400
transform 1 0 29344 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_254
timestamp 1669390400
transform 1 0 29792 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_266
timestamp 1669390400
transform 1 0 31136 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_276
timestamp 1669390400
transform 1 0 32256 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_284
timestamp 1669390400
transform 1 0 33152 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_291
timestamp 1669390400
transform 1 0 33936 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_295
timestamp 1669390400
transform 1 0 34384 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_299
timestamp 1669390400
transform 1 0 34832 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_303
timestamp 1669390400
transform 1 0 35280 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_307
timestamp 1669390400
transform 1 0 35728 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_311
timestamp 1669390400
transform 1 0 36176 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_315
timestamp 1669390400
transform 1 0 36624 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_321
timestamp 1669390400
transform 1 0 37296 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_324
timestamp 1669390400
transform 1 0 37632 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_328
timestamp 1669390400
transform 1 0 38080 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_332
timestamp 1669390400
transform 1 0 38528 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_336
timestamp 1669390400
transform 1 0 38976 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_368
timestamp 1669390400
transform 1 0 42560 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_384
timestamp 1669390400
transform 1 0 44352 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_388
timestamp 1669390400
transform 1 0 44800 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1669390400
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1669390400
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1669390400
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1669390400
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1669390400
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1669390400
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1669390400
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_598
timestamp 1669390400
transform 1 0 68320 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1669390400
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_605
timestamp 1669390400
transform 1 0 69104 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_669
timestamp 1669390400
transform 1 0 76272 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1669390400
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_676
timestamp 1669390400
transform 1 0 77056 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_684
timestamp 1669390400
transform 1 0 77952 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_6
timestamp 1669390400
transform 1 0 2016 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_10
timestamp 1669390400
transform 1 0 2464 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_14
timestamp 1669390400
transform 1 0 2912 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_18
timestamp 1669390400
transform 1 0 3360 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_22
timestamp 1669390400
transform 1 0 3808 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_30
timestamp 1669390400
transform 1 0 4704 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_40
timestamp 1669390400
transform 1 0 5824 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_50
timestamp 1669390400
transform 1 0 6944 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_60
timestamp 1669390400
transform 1 0 8064 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_70
timestamp 1669390400
transform 1 0 9184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_73
timestamp 1669390400
transform 1 0 9520 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_86
timestamp 1669390400
transform 1 0 10976 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_98
timestamp 1669390400
transform 1 0 12320 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_110
timestamp 1669390400
transform 1 0 13664 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1669390400
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_144
timestamp 1669390400
transform 1 0 17472 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_155
timestamp 1669390400
transform 1 0 18704 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_157
timestamp 1669390400
transform 1 0 18928 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_164
timestamp 1669390400
transform 1 0 19712 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_197
timestamp 1669390400
transform 1 0 23408 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_207
timestamp 1669390400
transform 1 0 24528 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_209
timestamp 1669390400
transform 1 0 24752 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1669390400
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_215
timestamp 1669390400
transform 1 0 25424 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_245
timestamp 1669390400
transform 1 0 28784 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_262
timestamp 1669390400
transform 1 0 30688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_279
timestamp 1669390400
transform 1 0 32592 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1669390400
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_286
timestamp 1669390400
transform 1 0 33376 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_299
timestamp 1669390400
transform 1 0 34832 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_303
timestamp 1669390400
transform 1 0 35280 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_307
timestamp 1669390400
transform 1 0 35728 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_311
timestamp 1669390400
transform 1 0 36176 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_315
timestamp 1669390400
transform 1 0 36624 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_319
timestamp 1669390400
transform 1 0 37072 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_323
timestamp 1669390400
transform 1 0 37520 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_327
timestamp 1669390400
transform 1 0 37968 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_331
timestamp 1669390400
transform 1 0 38416 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_335
timestamp 1669390400
transform 1 0 38864 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_339
timestamp 1669390400
transform 1 0 39312 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_343
timestamp 1669390400
transform 1 0 39760 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_351
timestamp 1669390400
transform 1 0 40656 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1669390400
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1669390400
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1669390400
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1669390400
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1669390400
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1669390400
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1669390400
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_570
timestamp 1669390400
transform 1 0 65184 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_634
timestamp 1669390400
transform 1 0 72352 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1669390400
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_641
timestamp 1669390400
transform 1 0 73136 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_673
timestamp 1669390400
transform 1 0 76720 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_681
timestamp 1669390400
transform 1 0 77616 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_685
timestamp 1669390400
transform 1 0 78064 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_687
timestamp 1669390400
transform 1 0 78288 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_8
timestamp 1669390400
transform 1 0 2240 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_12
timestamp 1669390400
transform 1 0 2688 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_16
timestamp 1669390400
transform 1 0 3136 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_20
timestamp 1669390400
transform 1 0 3584 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_24
timestamp 1669390400
transform 1 0 4032 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1669390400
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_37
timestamp 1669390400
transform 1 0 5488 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_47
timestamp 1669390400
transform 1 0 6608 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_61
timestamp 1669390400
transform 1 0 8176 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_63
timestamp 1669390400
transform 1 0 8400 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_70
timestamp 1669390400
transform 1 0 9184 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_80
timestamp 1669390400
transform 1 0 10304 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_97
timestamp 1669390400
transform 1 0 12208 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1669390400
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_108
timestamp 1669390400
transform 1 0 13440 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_138
timestamp 1669390400
transform 1 0 16800 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_169
timestamp 1669390400
transform 1 0 20272 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1669390400
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_179
timestamp 1669390400
transform 1 0 21392 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_189
timestamp 1669390400
transform 1 0 22512 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_193
timestamp 1669390400
transform 1 0 22960 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_226
timestamp 1669390400
transform 1 0 26656 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_244
timestamp 1669390400
transform 1 0 28672 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_250
timestamp 1669390400
transform 1 0 29344 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_266
timestamp 1669390400
transform 1 0 31136 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_270
timestamp 1669390400
transform 1 0 31584 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_306
timestamp 1669390400
transform 1 0 35616 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_310
timestamp 1669390400
transform 1 0 36064 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_314
timestamp 1669390400
transform 1 0 36512 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1669390400
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_321
timestamp 1669390400
transform 1 0 37296 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_324
timestamp 1669390400
transform 1 0 37632 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_328
timestamp 1669390400
transform 1 0 38080 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_332
timestamp 1669390400
transform 1 0 38528 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_336
timestamp 1669390400
transform 1 0 38976 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_340
timestamp 1669390400
transform 1 0 39424 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_344
timestamp 1669390400
transform 1 0 39872 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_348
timestamp 1669390400
transform 1 0 40320 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_380
timestamp 1669390400
transform 1 0 43904 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_388
timestamp 1669390400
transform 1 0 44800 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1669390400
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1669390400
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1669390400
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1669390400
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1669390400
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1669390400
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1669390400
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_605
timestamp 1669390400
transform 1 0 69104 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_669
timestamp 1669390400
transform 1 0 76272 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1669390400
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_676
timestamp 1669390400
transform 1 0 77056 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_684
timestamp 1669390400
transform 1 0 77952 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_6
timestamp 1669390400
transform 1 0 2016 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_10
timestamp 1669390400
transform 1 0 2464 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_18
timestamp 1669390400
transform 1 0 3360 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_51
timestamp 1669390400
transform 1 0 7056 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_53
timestamp 1669390400
transform 1 0 7280 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_60
timestamp 1669390400
transform 1 0 8064 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_70
timestamp 1669390400
transform 1 0 9184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_73
timestamp 1669390400
transform 1 0 9520 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_75
timestamp 1669390400
transform 1 0 9744 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_84
timestamp 1669390400
transform 1 0 10752 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_96
timestamp 1669390400
transform 1 0 12096 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_109
timestamp 1669390400
transform 1 0 13552 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_111
timestamp 1669390400
transform 1 0 13776 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1669390400
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_144
timestamp 1669390400
transform 1 0 17472 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_161
timestamp 1669390400
transform 1 0 19376 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_163
timestamp 1669390400
transform 1 0 19600 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_166
timestamp 1669390400
transform 1 0 19936 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_199
timestamp 1669390400
transform 1 0 23632 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1669390400
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_215
timestamp 1669390400
transform 1 0 25424 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_245
timestamp 1669390400
transform 1 0 28784 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_249
timestamp 1669390400
transform 1 0 29232 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1669390400
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_286
timestamp 1669390400
transform 1 0 33376 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_298
timestamp 1669390400
transform 1 0 34720 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_302
timestamp 1669390400
transform 1 0 35168 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_306
timestamp 1669390400
transform 1 0 35616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_310
timestamp 1669390400
transform 1 0 36064 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_314
timestamp 1669390400
transform 1 0 36512 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_318
timestamp 1669390400
transform 1 0 36960 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_322
timestamp 1669390400
transform 1 0 37408 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_326
timestamp 1669390400
transform 1 0 37856 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_330
timestamp 1669390400
transform 1 0 38304 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_334
timestamp 1669390400
transform 1 0 38752 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_338
timestamp 1669390400
transform 1 0 39200 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_342
timestamp 1669390400
transform 1 0 39648 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_346
timestamp 1669390400
transform 1 0 40096 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_350
timestamp 1669390400
transform 1 0 40544 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1669390400
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_357
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_360
timestamp 1669390400
transform 1 0 41664 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_424
timestamp 1669390400
transform 1 0 48832 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1669390400
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1669390400
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1669390400
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1669390400
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1669390400
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1669390400
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1669390400
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1669390400
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1669390400
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_641
timestamp 1669390400
transform 1 0 73136 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_673
timestamp 1669390400
transform 1 0 76720 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_681
timestamp 1669390400
transform 1 0 77616 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_685
timestamp 1669390400
transform 1 0 78064 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_687
timestamp 1669390400
transform 1 0 78288 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_4
timestamp 1669390400
transform 1 0 1792 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_15
timestamp 1669390400
transform 1 0 3024 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_21
timestamp 1669390400
transform 1 0 3696 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_34
timestamp 1669390400
transform 1 0 5152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_70
timestamp 1669390400
transform 1 0 9184 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_74
timestamp 1669390400
transform 1 0 9632 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1669390400
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_108
timestamp 1669390400
transform 1 0 13440 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_114
timestamp 1669390400
transform 1 0 14112 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_147
timestamp 1669390400
transform 1 0 17808 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_157
timestamp 1669390400
transform 1 0 18928 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_159
timestamp 1669390400
transform 1 0 19152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1669390400
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_179
timestamp 1669390400
transform 1 0 21392 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_183
timestamp 1669390400
transform 1 0 21840 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_214
timestamp 1669390400
transform 1 0 25312 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1669390400
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_250
timestamp 1669390400
transform 1 0 29344 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_256
timestamp 1669390400
transform 1 0 30016 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_270
timestamp 1669390400
transform 1 0 31584 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_304
timestamp 1669390400
transform 1 0 35392 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_312
timestamp 1669390400
transform 1 0 36288 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_316
timestamp 1669390400
transform 1 0 36736 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1669390400
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_321
timestamp 1669390400
transform 1 0 37296 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_324
timestamp 1669390400
transform 1 0 37632 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_328
timestamp 1669390400
transform 1 0 38080 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_332
timestamp 1669390400
transform 1 0 38528 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_336
timestamp 1669390400
transform 1 0 38976 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_340
timestamp 1669390400
transform 1 0 39424 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_344
timestamp 1669390400
transform 1 0 39872 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_348
timestamp 1669390400
transform 1 0 40320 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_352
timestamp 1669390400
transform 1 0 40768 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_356
timestamp 1669390400
transform 1 0 41216 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_360
timestamp 1669390400
transform 1 0 41664 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_364
timestamp 1669390400
transform 1 0 42112 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_380
timestamp 1669390400
transform 1 0 43904 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_388
timestamp 1669390400
transform 1 0 44800 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1669390400
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1669390400
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_463
timestamp 1669390400
transform 1 0 53200 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_471
timestamp 1669390400
transform 1 0 54096 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_475
timestamp 1669390400
transform 1 0 54544 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_477
timestamp 1669390400
transform 1 0 54768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_480
timestamp 1669390400
transform 1 0 55104 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_498
timestamp 1669390400
transform 1 0 57120 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_530
timestamp 1669390400
transform 1 0 60704 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1669390400
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1669390400
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1669390400
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_605
timestamp 1669390400
transform 1 0 69104 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_637
timestamp 1669390400
transform 1 0 72688 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_653
timestamp 1669390400
transform 1 0 74480 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_655
timestamp 1669390400
transform 1 0 74704 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_672
timestamp 1669390400
transform 1 0 76608 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_676
timestamp 1669390400
transform 1 0 77056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_679
timestamp 1669390400
transform 1 0 77392 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_687
timestamp 1669390400
transform 1 0 78288 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_4
timestamp 1669390400
transform 1 0 1792 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_7
timestamp 1669390400
transform 1 0 2128 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_11
timestamp 1669390400
transform 1 0 2576 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_15
timestamp 1669390400
transform 1 0 3024 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_23
timestamp 1669390400
transform 1 0 3920 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_33
timestamp 1669390400
transform 1 0 5040 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_37
timestamp 1669390400
transform 1 0 5488 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_41
timestamp 1669390400
transform 1 0 5936 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_51
timestamp 1669390400
transform 1 0 7056 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_69
timestamp 1669390400
transform 1 0 9072 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_72
timestamp 1669390400
transform 1 0 9408 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_86
timestamp 1669390400
transform 1 0 10976 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_104
timestamp 1669390400
transform 1 0 12992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_107
timestamp 1669390400
transform 1 0 13328 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_109
timestamp 1669390400
transform 1 0 13552 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_139
timestamp 1669390400
transform 1 0 16912 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_142
timestamp 1669390400
transform 1 0 17248 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_144
timestamp 1669390400
transform 1 0 17472 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_174
timestamp 1669390400
transform 1 0 20832 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_177
timestamp 1669390400
transform 1 0 21168 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_207
timestamp 1669390400
transform 1 0 24528 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_209
timestamp 1669390400
transform 1 0 24752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_212
timestamp 1669390400
transform 1 0 25088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_242
timestamp 1669390400
transform 1 0 28448 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_244
timestamp 1669390400
transform 1 0 28672 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_247
timestamp 1669390400
transform 1 0 29008 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_264
timestamp 1669390400
transform 1 0 30912 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_276
timestamp 1669390400
transform 1 0 32256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_282
timestamp 1669390400
transform 1 0 32928 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_285
timestamp 1669390400
transform 1 0 33264 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_303
timestamp 1669390400
transform 1 0 35280 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_307
timestamp 1669390400
transform 1 0 35728 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_311
timestamp 1669390400
transform 1 0 36176 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_317
timestamp 1669390400
transform 1 0 36848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_320
timestamp 1669390400
transform 1 0 37184 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_324
timestamp 1669390400
transform 1 0 37632 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_342
timestamp 1669390400
transform 1 0 39648 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_346
timestamp 1669390400
transform 1 0 40096 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_352
timestamp 1669390400
transform 1 0 40768 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_355
timestamp 1669390400
transform 1 0 41104 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_359
timestamp 1669390400
transform 1 0 41552 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_363
timestamp 1669390400
transform 1 0 42000 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_381
timestamp 1669390400
transform 1 0 44016 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_387
timestamp 1669390400
transform 1 0 44688 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_419
timestamp 1669390400
transform 1 0 48272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_422
timestamp 1669390400
transform 1 0 48608 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_425
timestamp 1669390400
transform 1 0 48944 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_433
timestamp 1669390400
transform 1 0 49840 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_437
timestamp 1669390400
transform 1 0 50288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_454
timestamp 1669390400
transform 1 0 52192 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_457
timestamp 1669390400
transform 1 0 52528 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_460
timestamp 1669390400
transform 1 0 52864 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_476
timestamp 1669390400
transform 1 0 54656 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_484
timestamp 1669390400
transform 1 0 55552 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_488
timestamp 1669390400
transform 1 0 56000 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_492
timestamp 1669390400
transform 1 0 56448 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_508
timestamp 1669390400
transform 1 0 58240 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_516
timestamp 1669390400
transform 1 0 59136 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_520
timestamp 1669390400
transform 1 0 59584 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_524
timestamp 1669390400
transform 1 0 60032 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_527
timestamp 1669390400
transform 1 0 60368 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_544
timestamp 1669390400
transform 1 0 62272 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_552
timestamp 1669390400
transform 1 0 63168 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_556
timestamp 1669390400
transform 1 0 63616 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_559
timestamp 1669390400
transform 1 0 63952 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_562
timestamp 1669390400
transform 1 0 64288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_579
timestamp 1669390400
transform 1 0 66192 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_587
timestamp 1669390400
transform 1 0 67088 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_591
timestamp 1669390400
transform 1 0 67536 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_594
timestamp 1669390400
transform 1 0 67872 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_597
timestamp 1669390400
transform 1 0 68208 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_615
timestamp 1669390400
transform 1 0 70224 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_623
timestamp 1669390400
transform 1 0 71120 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_627
timestamp 1669390400
transform 1 0 71568 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_629
timestamp 1669390400
transform 1 0 71792 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_632
timestamp 1669390400
transform 1 0 72128 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_636
timestamp 1669390400
transform 1 0 72576 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_654
timestamp 1669390400
transform 1 0 74592 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_662
timestamp 1669390400
transform 1 0 75488 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_664
timestamp 1669390400
transform 1 0 75712 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_667
timestamp 1669390400
transform 1 0 76048 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_683
timestamp 1669390400
transform 1 0 77840 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_687
timestamp 1669390400
transform 1 0 78288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1669390400
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1669390400
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1669390400
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1669390400
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1669390400
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1669390400
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1669390400
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1669390400
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1669390400
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1669390400
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1669390400
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1669390400
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1669390400
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1669390400
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1669390400
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1669390400
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1669390400
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1669390400
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1669390400
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1669390400
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1669390400
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1669390400
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1669390400
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1669390400
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1669390400
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1669390400
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1669390400
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1669390400
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1669390400
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1669390400
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1669390400
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1669390400
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1669390400
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1669390400
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1669390400
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1669390400
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1669390400
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1669390400
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1669390400
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1669390400
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1669390400
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1669390400
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1669390400
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1669390400
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1669390400
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1669390400
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1669390400
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1669390400
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1669390400
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1669390400
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1669390400
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1669390400
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1669390400
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1669390400
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1669390400
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1669390400
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1669390400
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1669390400
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1669390400
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1669390400
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1669390400
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1669390400
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1669390400
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1669390400
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1669390400
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1669390400
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1669390400
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1669390400
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1669390400
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1669390400
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1669390400
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1669390400
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1669390400
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1669390400
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1669390400
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1669390400
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1669390400
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1669390400
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1669390400
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1669390400
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1669390400
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1669390400
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1669390400
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1669390400
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1669390400
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1669390400
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1669390400
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1669390400
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1669390400
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1669390400
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1669390400
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1669390400
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1669390400
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1669390400
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1669390400
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1669390400
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1669390400
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1669390400
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1669390400
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1669390400
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1669390400
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1669390400
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1669390400
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1669390400
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1669390400
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1669390400
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1669390400
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1669390400
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1669390400
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1669390400
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1669390400
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1669390400
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1669390400
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1669390400
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1669390400
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1669390400
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1669390400
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1669390400
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1669390400
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1669390400
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1669390400
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1669390400
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1669390400
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1669390400
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1669390400
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1669390400
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1669390400
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1669390400
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1669390400
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1669390400
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1669390400
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1669390400
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1669390400
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1669390400
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1669390400
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1669390400
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1669390400
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1669390400
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1669390400
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1669390400
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1669390400
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1669390400
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1669390400
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1669390400
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1669390400
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1669390400
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1669390400
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1669390400
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1669390400
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1669390400
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1669390400
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1669390400
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1669390400
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1669390400
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1669390400
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1669390400
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1669390400
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1669390400
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1669390400
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1669390400
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1669390400
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1669390400
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1669390400
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1669390400
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1669390400
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1669390400
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1669390400
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1669390400
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1669390400
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1669390400
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1669390400
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1669390400
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1669390400
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1669390400
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1669390400
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1669390400
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1669390400
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1669390400
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1669390400
transform 1 0 5264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1669390400
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1669390400
transform 1 0 13104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1669390400
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1669390400
transform 1 0 20944 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1669390400
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1669390400
transform 1 0 28784 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1669390400
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1669390400
transform 1 0 36624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1669390400
transform 1 0 40544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1669390400
transform 1 0 44464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1669390400
transform 1 0 48384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1669390400
transform 1 0 52304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1669390400
transform 1 0 56224 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1669390400
transform 1 0 60144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1669390400
transform 1 0 64064 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1669390400
transform 1 0 67984 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1669390400
transform 1 0 71904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1669390400
transform 1 0 75824 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _246_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _247_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10864 0 -1 65856
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _248_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _249_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4592 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _250_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _251_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14672 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _252_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12096 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7840 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _254_
timestamp 1669390400
transform 1 0 10864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _255_
timestamp 1669390400
transform 1 0 11200 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _256_
timestamp 1669390400
transform 1 0 15008 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1669390400
transform 1 0 16128 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _258_
timestamp 1669390400
transform 1 0 18480 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _259_
timestamp 1669390400
transform 1 0 19488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _260_
timestamp 1669390400
transform 1 0 23072 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _261_
timestamp 1669390400
transform 1 0 24192 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _262_
timestamp 1669390400
transform 1 0 27664 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1669390400
transform 1 0 29120 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _264_
timestamp 1669390400
transform 1 0 32928 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _265_
timestamp 1669390400
transform 1 0 34160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _266_
timestamp 1669390400
transform 1 0 34608 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1669390400
transform 1 0 38192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _268_
timestamp 1669390400
transform 1 0 40320 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1669390400
transform 1 0 43344 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _270_
timestamp 1669390400
transform 1 0 47600 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _271_
timestamp 1669390400
transform 1 0 49392 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _272_
timestamp 1669390400
transform 1 0 52752 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _273_
timestamp 1669390400
transform 1 0 53872 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _274_
timestamp 1669390400
transform 1 0 52080 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _275_
timestamp 1669390400
transform 1 0 54768 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _276_
timestamp 1669390400
transform 1 0 51632 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1669390400
transform 1 0 57792 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _278_
timestamp 1669390400
transform 1 0 52640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _279_
timestamp 1669390400
transform 1 0 65744 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _280_
timestamp 1669390400
transform 1 0 17808 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1669390400
transform 1 0 29456 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _282_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8960 0 1 72128
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _283_
timestamp 1669390400
transform -1 0 28560 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _284_
timestamp 1669390400
transform 1 0 30128 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _285_
timestamp 1669390400
transform 1 0 6608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _286_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11536 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _287_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 9184 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _288_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3024 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _289_
timestamp 1669390400
transform 1 0 21952 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _290_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23072 0 1 67424
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _291_
timestamp 1669390400
transform -1 0 21056 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _292_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 30576 0 1 70560
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _293_
timestamp 1669390400
transform 1 0 17584 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _294_
timestamp 1669390400
transform -1 0 31136 0 1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _295_
timestamp 1669390400
transform -1 0 34720 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _296_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 25088 0 -1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _297_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10640 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _298_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22624 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _299_
timestamp 1669390400
transform -1 0 18704 0 -1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _300_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11536 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _301_
timestamp 1669390400
transform -1 0 6608 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _302_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13552 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _303_
timestamp 1669390400
transform -1 0 14672 0 1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _304_
timestamp 1669390400
transform 1 0 14784 0 -1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _305_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16464 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _306_
timestamp 1669390400
transform 1 0 21504 0 1 73696
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _307_
timestamp 1669390400
transform 1 0 21504 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _308_
timestamp 1669390400
transform 1 0 9632 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _309_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11200 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _310_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 13104 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _311_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11200 0 -1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _312_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9968 0 -1 73696
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _313_
timestamp 1669390400
transform -1 0 8960 0 -1 70560
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _314_
timestamp 1669390400
transform -1 0 7728 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _315_
timestamp 1669390400
transform -1 0 3920 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _316_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6832 0 1 70560
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _317_
timestamp 1669390400
transform -1 0 5824 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _318_
timestamp 1669390400
transform 1 0 5824 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _319_
timestamp 1669390400
transform 1 0 6720 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _320_
timestamp 1669390400
transform 1 0 8288 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _321_
timestamp 1669390400
transform 1 0 4256 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _322_
timestamp 1669390400
transform 1 0 9968 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _323_
timestamp 1669390400
transform -1 0 9184 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _324_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 2688 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _325_
timestamp 1669390400
transform -1 0 6048 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _326_
timestamp 1669390400
transform 1 0 13552 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _327_
timestamp 1669390400
transform 1 0 5264 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _328_
timestamp 1669390400
transform -1 0 13552 0 -1 75264
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _329_
timestamp 1669390400
transform -1 0 5040 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _330_
timestamp 1669390400
transform 1 0 7168 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _331_
timestamp 1669390400
transform 1 0 7504 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _332_
timestamp 1669390400
transform 1 0 10304 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _333_
timestamp 1669390400
transform -1 0 32256 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _334_
timestamp 1669390400
transform -1 0 8064 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _335_
timestamp 1669390400
transform 1 0 10640 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _336_
timestamp 1669390400
transform -1 0 19936 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _337_
timestamp 1669390400
transform -1 0 32256 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _338_
timestamp 1669390400
transform -1 0 18816 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _339_
timestamp 1669390400
transform -1 0 17136 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _340_
timestamp 1669390400
transform -1 0 10752 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _341_
timestamp 1669390400
transform 1 0 9408 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _342_
timestamp 1669390400
transform 1 0 8848 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _343_
timestamp 1669390400
transform -1 0 5152 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _344_
timestamp 1669390400
transform -1 0 28896 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _345_
timestamp 1669390400
transform 1 0 8288 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _346_
timestamp 1669390400
transform 1 0 10976 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _347_
timestamp 1669390400
transform -1 0 6608 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _348_
timestamp 1669390400
transform 1 0 18928 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _349_
timestamp 1669390400
transform 1 0 7952 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _350_
timestamp 1669390400
transform 1 0 5264 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _351_
timestamp 1669390400
transform -1 0 6944 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _352_
timestamp 1669390400
transform -1 0 10976 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _353_
timestamp 1669390400
transform 1 0 12208 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _354_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3136 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _355_
timestamp 1669390400
transform -1 0 8960 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _356_
timestamp 1669390400
transform 1 0 2912 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _357_
timestamp 1669390400
transform 1 0 9856 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _358_
timestamp 1669390400
transform 1 0 15568 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _359_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 18816 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _360_
timestamp 1669390400
transform -1 0 19824 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _361_
timestamp 1669390400
transform 1 0 27104 0 -1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _362_
timestamp 1669390400
transform 1 0 17920 0 1 72128
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _363_
timestamp 1669390400
transform 1 0 12208 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _364_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5824 0 1 64288
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _365_
timestamp 1669390400
transform 1 0 29456 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _366_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6832 0 1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _367_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1669390400
transform -1 0 5488 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _369_
timestamp 1669390400
transform 1 0 7280 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _370_
timestamp 1669390400
transform 1 0 6272 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _371_
timestamp 1669390400
transform 1 0 5824 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _372_
timestamp 1669390400
transform -1 0 7504 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _373_
timestamp 1669390400
transform 1 0 8624 0 1 68992
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _374_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11312 0 1 64288
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _375_
timestamp 1669390400
transform -1 0 5152 0 1 75264
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _376_
timestamp 1669390400
transform 1 0 4032 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _377_
timestamp 1669390400
transform -1 0 14112 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _378_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10976 0 1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _379_
timestamp 1669390400
transform 1 0 7168 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _380_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9296 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _381_
timestamp 1669390400
transform 1 0 9072 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _382_
timestamp 1669390400
transform -1 0 14896 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _383_
timestamp 1669390400
transform 1 0 2688 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _384_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12208 0 1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _385_
timestamp 1669390400
transform -1 0 9520 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _386_
timestamp 1669390400
transform 1 0 12992 0 -1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _387_
timestamp 1669390400
transform -1 0 13104 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _388_
timestamp 1669390400
transform 1 0 11872 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _389_
timestamp 1669390400
transform -1 0 12880 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _390_
timestamp 1669390400
transform 1 0 7952 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _391_
timestamp 1669390400
transform 1 0 13552 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _392_
timestamp 1669390400
transform -1 0 14112 0 -1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _393_
timestamp 1669390400
transform 1 0 10416 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _394_
timestamp 1669390400
transform -1 0 17136 0 1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _395_
timestamp 1669390400
transform 1 0 14784 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _396_
timestamp 1669390400
transform 1 0 13216 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _397_
timestamp 1669390400
transform -1 0 17024 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _398_
timestamp 1669390400
transform -1 0 15904 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _399_
timestamp 1669390400
transform 1 0 16576 0 1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _400_
timestamp 1669390400
transform -1 0 30128 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _401_
timestamp 1669390400
transform 1 0 26656 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _402_
timestamp 1669390400
transform -1 0 34384 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _403_
timestamp 1669390400
transform 1 0 25536 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _404_
timestamp 1669390400
transform 1 0 13552 0 1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _405_
timestamp 1669390400
transform 1 0 19488 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _406_
timestamp 1669390400
transform 1 0 18144 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _407_
timestamp 1669390400
transform 1 0 16240 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _408_
timestamp 1669390400
transform -1 0 11984 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _409_
timestamp 1669390400
transform 1 0 26544 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _410_
timestamp 1669390400
transform 1 0 25536 0 -1 68992
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _411_
timestamp 1669390400
transform -1 0 26432 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _412_
timestamp 1669390400
transform 1 0 12544 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _413_
timestamp 1669390400
transform -1 0 16352 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _414_
timestamp 1669390400
transform 1 0 17024 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _415_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17360 0 1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1669390400
transform 1 0 18368 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _417_
timestamp 1669390400
transform 1 0 20048 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _418_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20944 0 1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _419_
timestamp 1669390400
transform 1 0 21056 0 -1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _420_
timestamp 1669390400
transform 1 0 21728 0 1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _421_
timestamp 1669390400
transform -1 0 30688 0 -1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _422_
timestamp 1669390400
transform 1 0 23632 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _423_
timestamp 1669390400
transform 1 0 18032 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _424_
timestamp 1669390400
transform -1 0 22848 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _425_
timestamp 1669390400
transform -1 0 23184 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _426_
timestamp 1669390400
transform 1 0 24080 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _427_
timestamp 1669390400
transform 1 0 21840 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _428_
timestamp 1669390400
transform -1 0 20496 0 1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _429_
timestamp 1669390400
transform -1 0 13104 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _430_
timestamp 1669390400
transform -1 0 30016 0 -1 70560
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _431_
timestamp 1669390400
transform 1 0 17920 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _432_
timestamp 1669390400
transform -1 0 28672 0 1 64288
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _433_
timestamp 1669390400
transform 1 0 23744 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _434_
timestamp 1669390400
transform -1 0 26096 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _435_
timestamp 1669390400
transform -1 0 25424 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _436_
timestamp 1669390400
transform 1 0 24976 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _437_
timestamp 1669390400
transform 1 0 23072 0 -1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _438_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 28224 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1669390400
transform -1 0 19712 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _440_
timestamp 1669390400
transform -1 0 30016 0 -1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _441_
timestamp 1669390400
transform -1 0 30128 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _442_
timestamp 1669390400
transform -1 0 30800 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _443_
timestamp 1669390400
transform 1 0 26768 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _444_
timestamp 1669390400
transform 1 0 25536 0 -1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _445_
timestamp 1669390400
transform 1 0 27440 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _446_
timestamp 1669390400
transform -1 0 24528 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _447_
timestamp 1669390400
transform -1 0 24528 0 1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _448_
timestamp 1669390400
transform -1 0 26432 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _449_
timestamp 1669390400
transform 1 0 23296 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _450_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20720 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _451_
timestamp 1669390400
transform 1 0 26656 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _452_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26320 0 1 64288
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _453_
timestamp 1669390400
transform 1 0 27888 0 1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _454_
timestamp 1669390400
transform 1 0 31136 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _455_
timestamp 1669390400
transform -1 0 31808 0 1 65856
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _456_
timestamp 1669390400
transform -1 0 32032 0 -1 68992
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _457_
timestamp 1669390400
transform -1 0 26656 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _458_
timestamp 1669390400
transform 1 0 20160 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _459_
timestamp 1669390400
transform 1 0 30352 0 -1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _460_
timestamp 1669390400
transform 1 0 32256 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _461_
timestamp 1669390400
transform 1 0 31472 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _462_
timestamp 1669390400
transform -1 0 33040 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _463_
timestamp 1669390400
transform 1 0 30912 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _464_
timestamp 1669390400
transform 1 0 32032 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _465_
timestamp 1669390400
transform -1 0 33152 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _466_
timestamp 1669390400
transform 1 0 33488 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _467_
timestamp 1669390400
transform 1 0 32256 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _468_
timestamp 1669390400
transform 1 0 31920 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _469_
timestamp 1669390400
transform -1 0 33936 0 1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _470_
timestamp 1669390400
transform 1 0 30240 0 1 75264
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _471_
timestamp 1669390400
transform 1 0 31808 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _472_
timestamp 1669390400
transform -1 0 36288 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _473_
timestamp 1669390400
transform 1 0 29792 0 1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _474_
timestamp 1669390400
transform 1 0 33264 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _475_
timestamp 1669390400
transform 1 0 33488 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _476_
timestamp 1669390400
transform 1 0 32144 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _477_
timestamp 1669390400
transform 1 0 31136 0 -1 73696
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _478_
timestamp 1669390400
transform -1 0 33040 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _479_
timestamp 1669390400
transform 1 0 32480 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _480_
timestamp 1669390400
transform 1 0 26880 0 1 70560
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _481_
timestamp 1669390400
transform 1 0 33376 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _482_
timestamp 1669390400
transform 1 0 31584 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _483_
timestamp 1669390400
transform -1 0 30912 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _484_
timestamp 1669390400
transform 1 0 29008 0 -1 67424
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _485_
timestamp 1669390400
transform -1 0 30352 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _486_
timestamp 1669390400
transform -1 0 31024 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _487_
timestamp 1669390400
transform -1 0 29008 0 1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _488_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 28224 0 -1 68992
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _489_
timestamp 1669390400
transform 1 0 24304 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _490_
timestamp 1669390400
transform 1 0 21168 0 -1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _491_
timestamp 1669390400
transform -1 0 27552 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _492_
timestamp 1669390400
transform -1 0 27664 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _493_
timestamp 1669390400
transform -1 0 23072 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _494_
timestamp 1669390400
transform 1 0 11424 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _495_
timestamp 1669390400
transform -1 0 10752 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _496_
timestamp 1669390400
transform -1 0 11312 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _497_
timestamp 1669390400
transform 1 0 12544 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _498_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13104 0 -1 65856
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _499_
timestamp 1669390400
transform -1 0 17024 0 -1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _500_
timestamp 1669390400
transform -1 0 21056 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _501_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14896 0 1 67424
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _502_
timestamp 1669390400
transform -1 0 12320 0 1 65856
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _503_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 19152 0 -1 70560
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _504_
timestamp 1669390400
transform 1 0 7392 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _505_
timestamp 1669390400
transform -1 0 10752 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _506_
timestamp 1669390400
transform 1 0 7840 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _507_
timestamp 1669390400
transform 1 0 7728 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _508_
timestamp 1669390400
transform -1 0 8960 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1669390400
transform -1 0 7616 0 1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _510_
timestamp 1669390400
transform -1 0 7056 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _511_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 28448 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _512_
timestamp 1669390400
transform -1 0 28784 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _513_
timestamp 1669390400
transform -1 0 16800 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _514_
timestamp 1669390400
transform -1 0 28784 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _515_
timestamp 1669390400
transform -1 0 24752 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _516_
timestamp 1669390400
transform -1 0 24752 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _517_
timestamp 1669390400
transform 1 0 17024 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _518_
timestamp 1669390400
transform 1 0 17584 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _519_
timestamp 1669390400
transform 1 0 11312 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _520_
timestamp 1669390400
transform -1 0 17136 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _521_
timestamp 1669390400
transform -1 0 28784 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _522_
timestamp 1669390400
transform 1 0 13552 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _523_
timestamp 1669390400
transform 1 0 22064 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _524_
timestamp 1669390400
transform 1 0 9856 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _525_
timestamp 1669390400
transform 1 0 25088 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _526_
timestamp 1669390400
transform -1 0 20272 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _527_
timestamp 1669390400
transform -1 0 9184 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _528_
timestamp 1669390400
transform 1 0 22064 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _529_
timestamp 1669390400
transform -1 0 16800 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _530_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 29008 0 1 72128
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _531_
timestamp 1669390400
transform -1 0 24528 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _532_
timestamp 1669390400
transform 1 0 13328 0 -1 70560
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _533_
timestamp 1669390400
transform -1 0 21056 0 1 67424
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _534_
timestamp 1669390400
transform -1 0 23408 0 -1 70560
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _535_
timestamp 1669390400
transform 1 0 23184 0 1 73696
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _536_
timestamp 1669390400
transform 1 0 19152 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _537_
timestamp 1669390400
transform -1 0 9184 0 -1 68992
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _538_
timestamp 1669390400
transform -1 0 17808 0 1 75264
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _539_
timestamp 1669390400
transform 1 0 20160 0 -1 75264
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _540_
timestamp 1669390400
transform -1 0 17696 0 1 72128
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _541_
timestamp 1669390400
transform -1 0 11312 0 1 70560
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _542_
timestamp 1669390400
transform -1 0 16912 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _543_
timestamp 1669390400
transform -1 0 7056 0 -1 75264
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _544_
timestamp 1669390400
transform 1 0 19936 0 -1 73696
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _545_
timestamp 1669390400
transform 1 0 13888 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _546_
timestamp 1669390400
transform 1 0 9856 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _547_
timestamp 1669390400
transform -1 0 26544 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _548_
timestamp 1669390400
transform -1 0 29008 0 1 75264
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15120 0 1 70560
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform 1 0 19040 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform 1 0 19040 0 -1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform -1 0 52192 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 57120 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform -1 0 62272 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform -1 0 66192 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 70224 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform -1 0 74592 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform -1 0 12992 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform -1 0 19376 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform -1 0 21056 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 28672 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform -1 0 30912 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform -1 0 35280 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform -1 0 39648 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform -1 0 44016 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform -1 0 48272 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform -1 0 76608 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform 1 0 74816 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 3920 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform -1 0 50960 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 54096 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform 1 0 58464 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform 1 0 64400 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform 1 0 68320 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform 1 0 72912 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform 1 0 7056 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 11424 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 17360 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 21280 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 25872 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform 1 0 30576 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform 1 0 34944 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform 1 0 40880 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform 1 0 44800 0 1 3136
box -86 -86 1654 870
<< labels >>
flabel metal2 s 77504 0 77616 800 0 FreeSans 448 90 0 0 bs
port 0 nsew signal tristate
flabel metal2 s 2800 79200 2912 80000 0 FreeSans 448 90 0 0 clk
port 1 nsew signal input
flabel metal2 s 7168 79200 7280 80000 0 FreeSans 448 90 0 0 co[0]
port 2 nsew signal input
flabel metal2 s 50848 79200 50960 80000 0 FreeSans 448 90 0 0 co[10]
port 3 nsew signal input
flabel metal2 s 55216 79200 55328 80000 0 FreeSans 448 90 0 0 co[11]
port 4 nsew signal input
flabel metal2 s 59584 79200 59696 80000 0 FreeSans 448 90 0 0 co[12]
port 5 nsew signal input
flabel metal2 s 63952 79200 64064 80000 0 FreeSans 448 90 0 0 co[13]
port 6 nsew signal input
flabel metal2 s 68320 79200 68432 80000 0 FreeSans 448 90 0 0 co[14]
port 7 nsew signal input
flabel metal2 s 72688 79200 72800 80000 0 FreeSans 448 90 0 0 co[15]
port 8 nsew signal input
flabel metal2 s 11536 79200 11648 80000 0 FreeSans 448 90 0 0 co[1]
port 9 nsew signal input
flabel metal2 s 15904 79200 16016 80000 0 FreeSans 448 90 0 0 co[2]
port 10 nsew signal input
flabel metal2 s 20272 79200 20384 80000 0 FreeSans 448 90 0 0 co[3]
port 11 nsew signal input
flabel metal2 s 24640 79200 24752 80000 0 FreeSans 448 90 0 0 co[4]
port 12 nsew signal input
flabel metal2 s 29008 79200 29120 80000 0 FreeSans 448 90 0 0 co[5]
port 13 nsew signal input
flabel metal2 s 33376 79200 33488 80000 0 FreeSans 448 90 0 0 co[6]
port 14 nsew signal input
flabel metal2 s 37744 79200 37856 80000 0 FreeSans 448 90 0 0 co[7]
port 15 nsew signal input
flabel metal2 s 42112 79200 42224 80000 0 FreeSans 448 90 0 0 co[8]
port 16 nsew signal input
flabel metal2 s 46480 79200 46592 80000 0 FreeSans 448 90 0 0 co[9]
port 17 nsew signal input
flabel metal2 s 77056 79200 77168 80000 0 FreeSans 448 90 0 0 st
port 18 nsew signal input
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 20 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 20 nsew ground bidirectional
flabel metal2 s 2240 0 2352 800 0 FreeSans 448 90 0 0 x[0]
port 21 nsew signal tristate
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 x[10]
port 22 nsew signal tristate
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 x[11]
port 23 nsew signal tristate
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 x[12]
port 24 nsew signal tristate
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 x[13]
port 25 nsew signal tristate
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 x[14]
port 26 nsew signal tristate
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 x[15]
port 27 nsew signal tristate
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 x[1]
port 28 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 x[2]
port 29 nsew signal tristate
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 x[3]
port 30 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 x[4]
port 31 nsew signal tristate
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 x[5]
port 32 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 x[6]
port 33 nsew signal tristate
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 x[7]
port 34 nsew signal tristate
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 x[8]
port 35 nsew signal tristate
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 x[9]
port 36 nsew signal tristate
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 25368 73864 25368 73864 0 Datapath.i\[0\]
rlabel metal2 46872 5264 46872 5264 0 Datapath.i\[10\]
rlabel metal2 53368 5544 53368 5544 0 Datapath.i\[11\]
rlabel metal2 25144 76888 25144 76888 0 Datapath.i\[12\]
rlabel metal3 49336 4536 49336 4536 0 Datapath.i\[13\]
rlabel metal3 52248 3528 52248 3528 0 Datapath.i\[14\]
rlabel metal2 17192 65800 17192 65800 0 Datapath.i\[15\]
rlabel metal2 11928 4368 11928 4368 0 Datapath.i\[1\]
rlabel metal2 2632 60144 2632 60144 0 Datapath.i\[2\]
rlabel metal3 25648 74760 25648 74760 0 Datapath.i\[3\]
rlabel metal2 18648 5936 18648 5936 0 Datapath.i\[4\]
rlabel metal2 23016 5208 23016 5208 0 Datapath.i\[5\]
rlabel metal2 27552 4536 27552 4536 0 Datapath.i\[6\]
rlabel metal2 20664 76440 20664 76440 0 Datapath.i\[7\]
rlabel metal3 34552 5208 34552 5208 0 Datapath.i\[8\]
rlabel metal3 10528 48552 10528 48552 0 Datapath.i\[9\]
rlabel metal3 15512 61544 15512 61544 0 Datapath.k\[0\]
rlabel metal2 18200 75376 18200 75376 0 Datapath.k\[10\]
rlabel metal2 2688 73976 2688 73976 0 Datapath.k\[11\]
rlabel metal2 18088 66696 18088 66696 0 Datapath.k\[12\]
rlabel metal2 14504 72072 14504 72072 0 Datapath.k\[13\]
rlabel metal3 20160 74368 20160 74368 0 Datapath.k\[14\]
rlabel metal3 20160 76048 20160 76048 0 Datapath.k\[15\]
rlabel metal2 20888 69244 20888 69244 0 Datapath.k\[16\]
rlabel metal2 3192 63392 3192 63392 0 Datapath.k\[17\]
rlabel metal4 8568 72016 8568 72016 0 Datapath.k\[18\]
rlabel metal2 17640 70392 17640 70392 0 Datapath.k\[19\]
rlabel metal2 18704 74760 18704 74760 0 Datapath.k\[1\]
rlabel metal2 19880 58520 19880 58520 0 Datapath.k\[2\]
rlabel metal2 20440 71344 20440 71344 0 Datapath.k\[3\]
rlabel metal4 21448 64120 21448 64120 0 Datapath.k\[4\]
rlabel metal3 2632 64792 2632 64792 0 Datapath.k\[5\]
rlabel metal3 9912 68040 9912 68040 0 Datapath.k\[6\]
rlabel metal2 19768 74760 19768 74760 0 Datapath.k\[7\]
rlabel metal2 24304 62888 24304 62888 0 Datapath.k\[8\]
rlabel metal2 22288 66920 22288 66920 0 Datapath.k\[9\]
rlabel metal3 16296 63392 16296 63392 0 FSM.CS\[0\]
rlabel metal3 24416 75432 24416 75432 0 FSM.CS\[1\]
rlabel metal2 19208 65856 19208 65856 0 FSM.NS\[0\]
rlabel metal2 40152 76664 40152 76664 0 FSM.NS\[1\]
rlabel metal2 40936 77056 40936 77056 0 _000_
rlabel metal3 20160 77616 20160 77616 0 _001_
rlabel metal2 15848 65968 15848 65968 0 _002_
rlabel metal2 38808 74424 38808 74424 0 _003_
rlabel metal3 9184 73864 9184 73864 0 _004_
rlabel metal2 13832 72128 13832 72128 0 _005_
rlabel metal2 2184 75768 2184 75768 0 _006_
rlabel metal2 18144 58520 18144 58520 0 _007_
rlabel metal2 10920 61768 10920 61768 0 _008_
rlabel metal2 1960 72072 1960 72072 0 _009_
rlabel metal4 27720 54908 27720 54908 0 _010_
rlabel metal2 2408 77056 2408 77056 0 _011_
rlabel metal2 23016 77056 23016 77056 0 _012_
rlabel metal3 10416 72072 10416 72072 0 _013_
rlabel metal2 26040 68264 26040 68264 0 _014_
rlabel metal2 19096 75964 19096 75964 0 _015_
rlabel metal4 18200 61208 18200 61208 0 _016_
rlabel metal2 23016 69552 23016 69552 0 _017_
rlabel metal2 18312 63840 18312 63840 0 _018_
rlabel metal2 4200 73192 4200 73192 0 _019_
rlabel metal2 2520 77224 2520 77224 0 _020_
rlabel metal4 3192 65632 3192 65632 0 _021_
rlabel metal2 20104 68040 20104 68040 0 _022_
rlabel metal3 26152 69440 26152 69440 0 _023_
rlabel metal2 24080 73528 24080 73528 0 _024_
rlabel metal2 18144 71624 18144 71624 0 _025_
rlabel metal3 17976 65464 17976 65464 0 _026_
rlabel metal3 23128 75712 23128 75712 0 _027_
rlabel metal2 20776 74760 20776 74760 0 _028_
rlabel metal3 2240 71624 2240 71624 0 _029_
rlabel metal3 10472 70616 10472 70616 0 _030_
rlabel metal2 15960 76272 15960 76272 0 _031_
rlabel metal3 2184 74536 2184 74536 0 _032_
rlabel metal4 3080 55132 3080 55132 0 _033_
rlabel metal2 14840 73472 14840 73472 0 _034_
rlabel metal2 10808 69496 10808 69496 0 _035_
rlabel metal2 17976 69944 17976 69944 0 _036_
rlabel metal2 2352 60984 2352 60984 0 _037_
rlabel metal3 4984 62216 4984 62216 0 _038_
rlabel metal2 28056 4704 28056 4704 0 _039_
rlabel metal3 9520 4312 9520 4312 0 _040_
rlabel metal2 11536 5096 11536 5096 0 _041_
rlabel metal2 16016 4312 16016 4312 0 _042_
rlabel metal2 19600 4424 19600 4424 0 _043_
rlabel metal2 24080 4984 24080 4984 0 _044_
rlabel metal3 28840 4312 28840 4312 0 _045_
rlabel metal2 34272 4424 34272 4424 0 _046_
rlabel metal3 36848 4424 36848 4424 0 _047_
rlabel metal3 42280 4424 42280 4424 0 _048_
rlabel metal3 48944 4424 48944 4424 0 _049_
rlabel metal3 53760 4312 53760 4312 0 _050_
rlabel metal3 53872 4424 53872 4424 0 _051_
rlabel metal2 57960 4256 57960 4256 0 _052_
rlabel metal2 65352 3864 65352 3864 0 _053_
rlabel metal3 29232 55496 29232 55496 0 _054_
rlabel metal2 30688 60984 30688 60984 0 _055_
rlabel metal2 29848 61208 29848 61208 0 _056_
rlabel metal2 30408 60424 30408 60424 0 _057_
rlabel metal2 8848 67032 8848 67032 0 _058_
rlabel metal2 18424 74984 18424 74984 0 _059_
rlabel metal3 2464 75432 2464 75432 0 _060_
rlabel metal2 18032 72408 18032 72408 0 _061_
rlabel metal2 18480 74312 18480 74312 0 _062_
rlabel metal2 20944 73976 20944 73976 0 _063_
rlabel metal2 24248 74480 24248 74480 0 _064_
rlabel metal3 21504 73416 21504 73416 0 _065_
rlabel metal3 27552 74872 27552 74872 0 _066_
rlabel metal2 24920 75376 24920 75376 0 _067_
rlabel metal2 24920 74648 24920 74648 0 _068_
rlabel metal2 22288 73976 22288 73976 0 _069_
rlabel metal2 25144 72856 25144 72856 0 _070_
rlabel metal2 22120 74424 22120 74424 0 _071_
rlabel metal2 17192 66416 17192 66416 0 _072_
rlabel metal2 14336 70952 14336 70952 0 _073_
rlabel metal2 14504 67984 14504 67984 0 _074_
rlabel metal2 3080 77056 3080 77056 0 _075_
rlabel metal2 16128 66808 16128 66808 0 _076_
rlabel metal3 18704 61768 18704 61768 0 _077_
rlabel metal2 21896 64232 21896 64232 0 _078_
rlabel metal3 21084 62216 21084 62216 0 _079_
rlabel metal2 39032 74704 39032 74704 0 _080_
rlabel metal2 7168 70168 7168 70168 0 _081_
rlabel metal2 26152 72352 26152 72352 0 _082_
rlabel metal3 8008 70056 8008 70056 0 _083_
rlabel metal3 4872 75880 4872 75880 0 _084_
rlabel metal2 5936 72408 5936 72408 0 _085_
rlabel metal3 7504 72744 7504 72744 0 _086_
rlabel metal2 12600 73976 12600 73976 0 _087_
rlabel metal2 3192 61712 3192 61712 0 _088_
rlabel metal2 10248 69496 10248 69496 0 _089_
rlabel metal2 5208 70112 5208 70112 0 _090_
rlabel metal2 5768 69664 5768 69664 0 _091_
rlabel metal3 5152 76216 5152 76216 0 _092_
rlabel metal2 3304 61544 3304 61544 0 _093_
rlabel metal3 9072 67144 9072 67144 0 _094_
rlabel metal3 8064 72296 8064 72296 0 _095_
rlabel metal2 19768 72856 19768 72856 0 _096_
rlabel metal2 7672 64344 7672 64344 0 _097_
rlabel metal2 18368 68600 18368 68600 0 _098_
rlabel metal3 2856 63896 2856 63896 0 _099_
rlabel metal2 9744 73920 9744 73920 0 _100_
rlabel metal2 2576 61544 2576 61544 0 _101_
rlabel metal3 2296 61656 2296 61656 0 _102_
rlabel metal2 24584 76188 24584 76188 0 _103_
rlabel metal3 8512 72968 8512 72968 0 _104_
rlabel metal2 19096 64456 19096 64456 0 _105_
rlabel metal2 19208 64624 19208 64624 0 _106_
rlabel metal2 5432 65520 5432 65520 0 _107_
rlabel metal2 3416 68208 3416 68208 0 _108_
rlabel metal2 2408 67480 2408 67480 0 _109_
rlabel metal2 4200 71512 4200 71512 0 _110_
rlabel metal2 3192 65576 3192 65576 0 _111_
rlabel metal2 10136 61040 10136 61040 0 _112_
rlabel metal2 15848 62608 15848 62608 0 _113_
rlabel metal2 2856 69104 2856 69104 0 _114_
rlabel metal2 21784 75152 21784 75152 0 _115_
rlabel metal2 18424 71624 18424 71624 0 _116_
rlabel metal3 29064 63000 29064 63000 0 _117_
rlabel metal3 28308 61768 28308 61768 0 _118_
rlabel metal3 17696 63784 17696 63784 0 _119_
rlabel metal2 5208 68544 5208 68544 0 _120_
rlabel metal3 8624 66024 8624 66024 0 _121_
rlabel metal2 6664 66136 6664 66136 0 _122_
rlabel metal2 6888 67536 6888 67536 0 _123_
rlabel metal2 7224 68152 7224 68152 0 _124_
rlabel metal3 11536 69160 11536 69160 0 _125_
rlabel metal4 2632 66640 2632 66640 0 _126_
rlabel metal2 4200 74088 4200 74088 0 _127_
rlabel metal2 3248 74872 3248 74872 0 _128_
rlabel metal3 15008 63112 15008 63112 0 _129_
rlabel metal2 9800 64456 9800 64456 0 _130_
rlabel metal2 16576 62328 16576 62328 0 _131_
rlabel metal2 13832 62636 13832 62636 0 _132_
rlabel metal3 2240 74648 2240 74648 0 _133_
rlabel metal2 3248 69832 3248 69832 0 _134_
rlabel metal2 9352 66528 9352 66528 0 _135_
rlabel metal2 15736 64344 15736 64344 0 _136_
rlabel metal3 14056 63896 14056 63896 0 _137_
rlabel metal2 11984 64120 11984 64120 0 _138_
rlabel metal3 2996 66360 2996 66360 0 _139_
rlabel metal3 9464 62552 9464 62552 0 _140_
rlabel metal2 13832 61768 13832 61768 0 _141_
rlabel metal3 12432 62328 12432 62328 0 _142_
rlabel metal2 18536 63896 18536 63896 0 _143_
rlabel metal3 17192 62552 17192 62552 0 _144_
rlabel metal3 17192 61992 17192 61992 0 _145_
rlabel metal2 16464 62552 16464 62552 0 _146_
rlabel metal2 16856 64400 16856 64400 0 _147_
rlabel metal2 17808 64792 17808 64792 0 _148_
rlabel metal2 25592 69160 25592 69160 0 _149_
rlabel metal3 26656 71736 26656 71736 0 _150_
rlabel metal2 26376 71792 26376 71792 0 _151_
rlabel metal2 11480 68040 11480 68040 0 _152_
rlabel metal3 19656 64120 19656 64120 0 _153_
rlabel metal2 16408 64792 16408 64792 0 _154_
rlabel metal2 16520 64568 16520 64568 0 _155_
rlabel metal2 26040 69104 26040 69104 0 _156_
rlabel metal2 26824 65016 26824 65016 0 _157_
rlabel metal2 25928 68824 25928 68824 0 _158_
rlabel metal2 39144 70000 39144 70000 0 _159_
rlabel metal3 16464 64904 16464 64904 0 _160_
rlabel metal2 20328 65800 20328 65800 0 _161_
rlabel metal2 19880 64568 19880 64568 0 _162_
rlabel metal3 19544 64008 19544 64008 0 _163_
rlabel metal2 20552 64456 20552 64456 0 _164_
rlabel metal2 22232 64288 22232 64288 0 _165_
rlabel metal2 23464 65744 23464 65744 0 _166_
rlabel metal2 22904 68488 22904 68488 0 _167_
rlabel metal2 24360 73024 24360 73024 0 _168_
rlabel metal2 18256 71960 18256 71960 0 _169_
rlabel metal2 21672 67648 21672 67648 0 _170_
rlabel metal3 22456 63336 22456 63336 0 _171_
rlabel metal2 24360 63896 24360 63896 0 _172_
rlabel metal2 22120 65576 22120 65576 0 _173_
rlabel metal2 15064 69384 15064 69384 0 _174_
rlabel metal3 17136 71960 17136 71960 0 _175_
rlabel metal2 18760 71680 18760 71680 0 _176_
rlabel metal2 23912 65296 23912 65296 0 _177_
rlabel metal3 24696 63672 24696 63672 0 _178_
rlabel metal2 25256 63504 25256 63504 0 _179_
rlabel metal3 25928 64680 25928 64680 0 _180_
rlabel metal3 25592 64568 25592 64568 0 _181_
rlabel metal2 24360 68376 24360 68376 0 _182_
rlabel metal2 3304 72800 3304 72800 0 _183_
rlabel metal3 25144 65464 25144 65464 0 _184_
rlabel metal3 28392 66248 28392 66248 0 _185_
rlabel metal2 28168 65800 28168 65800 0 _186_
rlabel metal2 27048 65744 27048 65744 0 _187_
rlabel metal2 26712 65464 26712 65464 0 _188_
rlabel metal2 26040 66528 26040 66528 0 _189_
rlabel metal2 26264 67200 26264 67200 0 _190_
rlabel metal3 24864 64792 24864 64792 0 _191_
rlabel metal3 22512 65240 22512 65240 0 _192_
rlabel metal2 20216 65688 20216 65688 0 _193_
rlabel metal2 28280 66696 28280 66696 0 _194_
rlabel metal3 27720 64904 27720 64904 0 _195_
rlabel metal3 30464 67032 30464 67032 0 _196_
rlabel metal2 31640 68656 31640 68656 0 _197_
rlabel metal3 32032 68488 32032 68488 0 _198_
rlabel metal2 20216 76552 20216 76552 0 _199_
rlabel metal2 20888 71792 20888 71792 0 _200_
rlabel via2 31528 68600 31528 68600 0 _201_
rlabel metal2 32760 68488 32760 68488 0 _202_
rlabel metal2 31752 68488 31752 68488 0 _203_
rlabel metal3 32312 69608 32312 69608 0 _204_
rlabel metal2 32088 71176 32088 71176 0 _205_
rlabel metal2 32984 71232 32984 71232 0 _206_
rlabel metal3 33768 69384 33768 69384 0 _207_
rlabel metal2 33880 69496 33880 69496 0 _208_
rlabel metal2 33656 70952 33656 70952 0 _209_
rlabel metal3 32256 70952 32256 70952 0 _210_
rlabel metal2 31416 75600 31416 75600 0 _211_
rlabel metal3 34552 75544 34552 75544 0 _212_
rlabel metal3 32536 73304 32536 73304 0 _213_
rlabel metal3 33824 69608 33824 69608 0 _214_
rlabel metal3 33320 70392 33320 70392 0 _215_
rlabel metal3 32088 71960 32088 71960 0 _216_
rlabel metal2 32536 74648 32536 74648 0 _217_
rlabel metal2 32648 72632 32648 72632 0 _218_
rlabel metal2 28112 69608 28112 69608 0 _219_
rlabel metal2 31752 70168 31752 70168 0 _220_
rlabel metal2 30072 68880 30072 68880 0 _221_
rlabel metal2 30576 67032 30576 67032 0 _222_
rlabel metal2 29064 68992 29064 68992 0 _223_
rlabel metal3 30464 69272 30464 69272 0 _224_
rlabel metal2 29960 68656 29960 68656 0 _225_
rlabel metal3 27608 69384 27608 69384 0 _226_
rlabel metal2 24472 68152 24472 68152 0 _227_
rlabel metal2 24808 67872 24808 67872 0 _228_
rlabel metal2 21672 66528 21672 66528 0 _229_
rlabel metal2 27272 68880 27272 68880 0 _230_
rlabel metal2 22680 65968 22680 65968 0 _231_
rlabel metal2 16408 66976 16408 66976 0 _232_
rlabel metal2 10472 66248 10472 66248 0 _233_
rlabel metal3 12040 66024 12040 66024 0 _234_
rlabel metal3 13944 65464 13944 65464 0 _235_
rlabel metal3 16128 65464 16128 65464 0 _236_
rlabel metal2 16632 68432 16632 68432 0 _237_
rlabel metal2 15736 66976 15736 66976 0 _238_
rlabel metal2 18200 69888 18200 69888 0 _239_
rlabel metal3 11928 43624 11928 43624 0 _240_
rlabel metal3 9184 63224 9184 63224 0 _241_
rlabel metal2 8568 67816 8568 67816 0 _242_
rlabel metal2 8008 69832 8008 69832 0 _243_
rlabel metal2 6720 75880 6720 75880 0 _244_
rlabel metal3 6832 76440 6832 76440 0 _245_
rlabel metal2 77560 2478 77560 2478 0 bs
rlabel metal2 2464 79240 2464 79240 0 clk
rlabel metal2 19208 69720 19208 69720 0 clknet_0_clk
rlabel metal2 1904 74760 1904 74760 0 clknet_2_0__leaf_clk
rlabel metal2 16968 75264 16968 75264 0 clknet_2_1__leaf_clk
rlabel metal2 16520 68376 16520 68376 0 clknet_2_2__leaf_clk
rlabel metal2 22344 76048 22344 76048 0 clknet_2_3__leaf_clk
rlabel metal3 3920 64008 3920 64008 0 co[0]
rlabel metal3 51240 76552 51240 76552 0 co[10]
rlabel metal2 55160 75768 55160 75768 0 co[11]
rlabel metal2 59808 76664 59808 76664 0 co[12]
rlabel metal2 63952 76664 63952 76664 0 co[13]
rlabel metal2 67816 76720 67816 76720 0 co[14]
rlabel metal2 72632 76664 72632 76664 0 co[15]
rlabel metal2 16296 58576 16296 58576 0 co[1]
rlabel metal2 2072 77728 2072 77728 0 co[2]
rlabel metal2 2968 77616 2968 77616 0 co[3]
rlabel metal2 24696 77154 24696 77154 0 co[4]
rlabel metal2 39256 75376 39256 75376 0 co[5]
rlabel metal3 34048 76552 34048 76552 0 co[6]
rlabel metal2 37688 76664 37688 76664 0 co[7]
rlabel metal2 42056 76664 42056 76664 0 co[8]
rlabel metal3 47096 76552 47096 76552 0 co[9]
rlabel metal2 22120 62496 22120 62496 0 net1
rlabel metal2 2856 57736 2856 57736 0 net10
rlabel metal3 20160 74928 20160 74928 0 net11
rlabel metal3 30072 60984 30072 60984 0 net12
rlabel metal2 30184 71232 30184 71232 0 net13
rlabel metal2 25704 69104 25704 69104 0 net14
rlabel metal2 42392 75040 42392 75040 0 net15
rlabel metal2 46648 74368 46648 74368 0 net16
rlabel metal2 74984 76552 74984 76552 0 net17
rlabel metal3 76328 4312 76328 4312 0 net18
rlabel metal3 2352 3528 2352 3528 0 net19
rlabel metal2 50456 74088 50456 74088 0 net2
rlabel metal3 50232 4424 50232 4424 0 net20
rlabel metal2 54376 3976 54376 3976 0 net21
rlabel metal3 55356 4424 55356 4424 0 net22
rlabel metal3 61432 4424 61432 4424 0 net23
rlabel metal2 68488 3976 68488 3976 0 net24
rlabel metal3 75320 3528 75320 3528 0 net25
rlabel metal2 7336 3976 7336 3976 0 net26
rlabel metal2 11648 4872 11648 4872 0 net27
rlabel metal3 17080 4424 17080 4424 0 net28
rlabel metal2 21448 3976 21448 3976 0 net29
rlabel metal2 55384 74312 55384 74312 0 net3
rlabel metal3 25368 4872 25368 4872 0 net30
rlabel metal3 30184 4424 30184 4424 0 net31
rlabel metal2 34664 3976 34664 3976 0 net32
rlabel metal2 38696 3976 38696 3976 0 net33
rlabel metal2 43848 3976 43848 3976 0 net34
rlabel metal2 60648 75488 60648 75488 0 net4
rlabel metal2 64568 75208 64568 75208 0 net5
rlabel metal2 68600 76272 68600 76272 0 net6
rlabel metal2 72968 76496 72968 76496 0 net7
rlabel metal2 2632 74872 2632 74872 0 net8
rlabel metal2 17752 74928 17752 74928 0 net9
rlabel metal2 77168 75768 77168 75768 0 st
rlabel metal2 2296 2086 2296 2086 0 x[0]
rlabel metal2 49336 2086 49336 2086 0 x[10]
rlabel metal2 54040 2198 54040 2198 0 x[11]
rlabel metal2 58744 2198 58744 2198 0 x[12]
rlabel metal2 63448 2198 63448 2198 0 x[13]
rlabel metal2 68152 2198 68152 2198 0 x[14]
rlabel metal2 72856 2198 72856 2198 0 x[15]
rlabel metal2 7000 2198 7000 2198 0 x[1]
rlabel metal2 11704 2198 11704 2198 0 x[2]
rlabel metal2 16408 2198 16408 2198 0 x[3]
rlabel metal2 21112 2198 21112 2198 0 x[4]
rlabel metal2 25816 2198 25816 2198 0 x[5]
rlabel metal2 30520 2198 30520 2198 0 x[6]
rlabel metal2 35224 2198 35224 2198 0 x[7]
rlabel metal2 39928 2198 39928 2198 0 x[8]
rlabel metal2 44632 2030 44632 2030 0 x[9]
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
