magic
tech gf180mcuC
magscale 1 5
timestamp 1670102150
<< obsm1 >>
rect 672 1538 39312 38849
<< metal2 >>
rect 1400 39600 1456 40000
rect 3584 39600 3640 40000
rect 5768 39600 5824 40000
rect 7952 39600 8008 40000
rect 10136 39600 10192 40000
rect 12320 39600 12376 40000
rect 14504 39600 14560 40000
rect 16688 39600 16744 40000
rect 18872 39600 18928 40000
rect 21056 39600 21112 40000
rect 23240 39600 23296 40000
rect 25424 39600 25480 40000
rect 27608 39600 27664 40000
rect 29792 39600 29848 40000
rect 31976 39600 32032 40000
rect 34160 39600 34216 40000
rect 36344 39600 36400 40000
rect 38528 39600 38584 40000
rect 1120 0 1176 400
rect 3472 0 3528 400
rect 5824 0 5880 400
rect 8176 0 8232 400
rect 10528 0 10584 400
rect 12880 0 12936 400
rect 15232 0 15288 400
rect 17584 0 17640 400
rect 19936 0 19992 400
rect 22288 0 22344 400
rect 24640 0 24696 400
rect 26992 0 27048 400
rect 29344 0 29400 400
rect 31696 0 31752 400
rect 34048 0 34104 400
rect 36400 0 36456 400
rect 38752 0 38808 400
<< obsm2 >>
rect 798 39570 1370 39975
rect 1486 39570 3554 39975
rect 3670 39570 5738 39975
rect 5854 39570 7922 39975
rect 8038 39570 10106 39975
rect 10222 39570 12290 39975
rect 12406 39570 14474 39975
rect 14590 39570 16658 39975
rect 16774 39570 18842 39975
rect 18958 39570 21026 39975
rect 21142 39570 23210 39975
rect 23326 39570 25394 39975
rect 25510 39570 27578 39975
rect 27694 39570 29762 39975
rect 29878 39570 31946 39975
rect 32062 39570 34130 39975
rect 34246 39570 36314 39975
rect 36430 39570 38498 39975
rect 38614 39570 38794 39975
rect 798 430 38794 39570
rect 798 400 1090 430
rect 1206 400 3442 430
rect 3558 400 5794 430
rect 5910 400 8146 430
rect 8262 400 10498 430
rect 10614 400 12850 430
rect 12966 400 15202 430
rect 15318 400 17554 430
rect 17670 400 19906 430
rect 20022 400 22258 430
rect 22374 400 24610 430
rect 24726 400 26962 430
rect 27078 400 29314 430
rect 29430 400 31666 430
rect 31782 400 34018 430
rect 34134 400 36370 430
rect 36486 400 38722 430
<< obsm3 >>
rect 569 1554 38799 39970
<< metal4 >>
rect 2224 1538 2384 38446
rect 9904 1538 10064 38446
rect 17584 1538 17744 38446
rect 25264 1538 25424 38446
rect 32944 1538 33104 38446
<< obsm4 >>
rect 574 38476 16842 39639
rect 574 1745 2194 38476
rect 2414 1745 9874 38476
rect 10094 1745 16842 38476
<< labels >>
rlabel metal2 s 38752 0 38808 400 6 bs
port 1 nsew signal output
rlabel metal2 s 1400 39600 1456 40000 6 clk
port 2 nsew signal input
rlabel metal2 s 3584 39600 3640 40000 6 co[0]
port 3 nsew signal input
rlabel metal2 s 25424 39600 25480 40000 6 co[10]
port 4 nsew signal input
rlabel metal2 s 27608 39600 27664 40000 6 co[11]
port 5 nsew signal input
rlabel metal2 s 29792 39600 29848 40000 6 co[12]
port 6 nsew signal input
rlabel metal2 s 31976 39600 32032 40000 6 co[13]
port 7 nsew signal input
rlabel metal2 s 34160 39600 34216 40000 6 co[14]
port 8 nsew signal input
rlabel metal2 s 36344 39600 36400 40000 6 co[15]
port 9 nsew signal input
rlabel metal2 s 5768 39600 5824 40000 6 co[1]
port 10 nsew signal input
rlabel metal2 s 7952 39600 8008 40000 6 co[2]
port 11 nsew signal input
rlabel metal2 s 10136 39600 10192 40000 6 co[3]
port 12 nsew signal input
rlabel metal2 s 12320 39600 12376 40000 6 co[4]
port 13 nsew signal input
rlabel metal2 s 14504 39600 14560 40000 6 co[5]
port 14 nsew signal input
rlabel metal2 s 16688 39600 16744 40000 6 co[6]
port 15 nsew signal input
rlabel metal2 s 18872 39600 18928 40000 6 co[7]
port 16 nsew signal input
rlabel metal2 s 21056 39600 21112 40000 6 co[8]
port 17 nsew signal input
rlabel metal2 s 23240 39600 23296 40000 6 co[9]
port 18 nsew signal input
rlabel metal2 s 38528 39600 38584 40000 6 st
port 19 nsew signal input
rlabel metal4 s 2224 1538 2384 38446 6 vdd
port 20 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 38446 6 vdd
port 20 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 38446 6 vdd
port 20 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 38446 6 vss
port 21 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 38446 6 vss
port 21 nsew ground bidirectional
rlabel metal2 s 1120 0 1176 400 6 x[0]
port 22 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 x[10]
port 23 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 x[11]
port 24 nsew signal output
rlabel metal2 s 29344 0 29400 400 6 x[12]
port 25 nsew signal output
rlabel metal2 s 31696 0 31752 400 6 x[13]
port 26 nsew signal output
rlabel metal2 s 34048 0 34104 400 6 x[14]
port 27 nsew signal output
rlabel metal2 s 36400 0 36456 400 6 x[15]
port 28 nsew signal output
rlabel metal2 s 3472 0 3528 400 6 x[1]
port 29 nsew signal output
rlabel metal2 s 5824 0 5880 400 6 x[2]
port 30 nsew signal output
rlabel metal2 s 8176 0 8232 400 6 x[3]
port 31 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 x[4]
port 32 nsew signal output
rlabel metal2 s 12880 0 12936 400 6 x[5]
port 33 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 x[6]
port 34 nsew signal output
rlabel metal2 s 17584 0 17640 400 6 x[7]
port 35 nsew signal output
rlabel metal2 s 19936 0 19992 400 6 x[8]
port 36 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 x[9]
port 37 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1652228
string GDS_FILE /home/dbarrios/collatz_wrap/openlane/collatz/runs/22_12_03_16_14/results/signoff/collatz.magic.gds
string GDS_START 239650
<< end >>

