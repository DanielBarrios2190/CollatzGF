* NGSPICE file created from collatz.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

.subckt collatz bs clk co[0] co[10] co[11] co[12] co[13] co[14] co[15] co[1] co[2]
+ co[3] co[4] co[5] co[6] co[7] co[8] co[9] st vdd vss x[0] x[10] x[11] x[12] x[13]
+ x[14] x[15] x[1] x[2] x[3] x[4] x[5] x[6] x[7] x[8] x[9]
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__429__I _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_501_ _042_ _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_432_ _040_ _037_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_363_ _047_ Datapath.i\[5\] _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__568__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__559__A1 _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_346_ _037_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_415_ Datapath.k\[14\] _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_680_ _315_ _311_ _320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__392__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__717__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_732_ _025_ clknet_2_2__leaf_clk Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_594_ _080_ _075_ _241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_663_ _222_ _303_ _304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput31 net31 x[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput20 net20 x[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_715_ _008_ clknet_2_0__leaf_clk Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__595__A2 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__347__A2 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_577_ _222_ _225_ _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_646_ Datapath.k\[15\] _103_ _038_ net6 _046_ _289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__360__I _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_500_ _103_ Datapath.k\[1\] _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_362_ _048_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_431_ _074_ _104_ FSM.NS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_629_ _270_ _272_ _273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__559__A2 _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_345_ FSM.CS\[1\] _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_414_ Datapath.k\[15\] _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__698__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__698__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__699__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__453__I _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__689__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__540__B1 _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_731_ _024_ clknet_2_2__leaf_clk Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_662_ _302_ _238_ _255_ _303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_593_ _221_ _238_ _239_ _240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I co[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__589__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput32 net32 x[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput21 net21 x[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_645_ _286_ _064_ _287_ _288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_714_ _007_ clknet_2_0__leaf_clk Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_576_ _223_ _224_ _225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__504__B1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I co[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__707__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__510__A3 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_361_ _047_ Datapath.i\[4\] _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_430_ _092_ _101_ _103_ _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_628_ _100_ _271_ _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_559_ _094_ _205_ _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__371__I Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_413_ Datapath.k\[5\] Datapath.k\[4\] _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_344_ FSM.CS\[0\] _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__477__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__468__A2 _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__395__A1 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__386__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__622__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__689__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__740__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__368__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__540__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_730_ _023_ clknet_2_2__leaf_clk Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_592_ _224_ _232_ _239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_661_ _301_ _302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__522__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__513__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput22 net22 x[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 x[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_713_ _006_ clknet_2_1__leaf_clk Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_644_ _278_ _280_ _284_ _287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_575_ Datapath.k\[8\] Datapath.k\[7\] _224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__504__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__369__I Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_360_ _046_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_558_ _204_ _207_ _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_627_ Datapath.k\[13\] Datapath.k\[12\] _271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_489_ _141_ Datapath.i\[13\] Datapath.i\[12\] Datapath.i\[11\] _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_412_ Datapath.k\[0\] _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__631__A3 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__395__A2 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__386__A2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__368__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_591_ _225_ _233_ _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_660_ _277_ _300_ _301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__390__I Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__522__A2 _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__589__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__513__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput34 net34 x[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 x[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__730__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_712_ _005_ clknet_2_1__leaf_clk Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_643_ _281_ _285_ _286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_574_ _076_ _213_ _223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__504__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__498__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__670__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_488_ _056_ _145_ _148_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_557_ _206_ _093_ _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_626_ _261_ _262_ _269_ _270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__489__A1 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__413__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_411_ _077_ _078_ _081_ _084_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_609_ _253_ _254_ _079_ _047_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_590_ _236_ _237_ _075_ _158_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 x[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_642_ _284_ _285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_711_ _004_ clknet_2_1__leaf_clk Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_573_ _221_ _222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_16_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__670__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__486__I _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_625_ _263_ _269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_556_ _205_ _206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_487_ _147_ _062_ _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I co[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__413__A2 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__720__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_410_ _082_ _083_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_608_ Datapath.k\[12\] _103_ _038_ net3 _046_ _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__743__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_539_ net12 _120_ Datapath.k\[6\] _102_ _042_ _191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__398__A1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__570__A1 _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__543__A1 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__525__A1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__516__A1 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__507__A1 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__530__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 x[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_641_ _282_ _283_ _284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_572_ _217_ _220_ _221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_710_ _003_ clknet_2_1__leaf_clk Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__541__B _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_555_ Datapath.k\[7\] Datapath.k\[6\] _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_624_ _267_ _268_ _099_ _047_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_486_ _146_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__646__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_538_ _185_ _188_ _189_ _190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_607_ _251_ _252_ _253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_469_ _131_ _053_ _062_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__398__A2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__570__A2 _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__561__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__710__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__623__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__733__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__470__A1 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__525__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__516__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__507__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 x[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_571_ _218_ _192_ _219_ _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_640_ Datapath.k\[14\] Datapath.k\[13\] _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__407__A1 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_485_ _143_ _056_ _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_554_ _200_ _195_ _204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_623_ Datapath.k\[13\] _103_ _038_ net4 _046_ _268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_8_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__646__B2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__646__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__489__A4 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__582__B1 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__628__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_468_ _052_ _129_ _132_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_537_ _185_ _188_ _060_ _189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_606_ _244_ _242_ _249_ _252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__564__B1 _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_399_ _060_ _037_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__398__A3 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__519__B1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__470__A2 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__691__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__443__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__723__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 x[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__539__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__434__A2 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_570_ _195_ _205_ _219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__370__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_699_ _336_ _337_ _121_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__361__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_622_ _264_ _064_ _266_ _267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_553_ _201_ _202_ _203_ _158_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_484_ _141_ Datapath.i\[11\] _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__646__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__582__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_605_ _250_ _036_ _251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__564__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_467_ _131_ _062_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_398_ _070_ _060_ net1 _071_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_536_ _187_ _087_ _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__555__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__546__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__537__A1 _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_519_ net10 _121_ Datapath.k\[4\] _102_ _042_ _173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__528__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__402__I Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__519__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__600__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput28 net28 x[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__571__B _219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_698_ _042_ Datapath.k\[18\] Datapath.k\[19\] _060_ _337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__361__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__391__B _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__655__A3 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_621_ _260_ _265_ _266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__591__A2 _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_483_ _055_ _140_ _144_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_552_ Datapath.k\[6\] _203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__713__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__405__I Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__736__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_535_ _186_ _184_ _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_604_ _244_ _242_ _249_ _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_466_ _128_ Datapath.i\[8\] Datapath.i\[7\] _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_397_ net8 net9 net10 net11 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__555__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__546__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__482__A1 _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_518_ _169_ _064_ _171_ _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__537__A2 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_449_ _117_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__473__A1 Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__528__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__464__A1 _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__519__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__437__B2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__479__B _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__600__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 bs vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net29 x[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__419__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__408__I Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__658__A1 _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_697_ _334_ _317_ _335_ _336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__656__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_551_ net13 _120_ Datapath.k\[7\] _102_ _046_ _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_620_ _262_ _263_ _265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_482_ _143_ _062_ _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__421__I Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_534_ Datapath.k\[5\] _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_465_ _051_ _127_ _130_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_603_ _081_ _248_ _249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_396_ _069_ net5 net6 net7 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_4_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__491__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__482__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_517_ _165_ _162_ _170_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_448_ _115_ Datapath.i\[4\] _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_379_ Datapath.i\[13\] _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__473__A2 Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__726__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__464__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__391__A1 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__382__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__373__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__600__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 x[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__419__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__355__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_696_ _329_ _333_ _335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__585__A1 _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_481_ _142_ Datapath.i\[11\] Datapath.i\[10\] _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_550_ _199_ _200_ _036_ _201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__567__A1 _214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_679_ _318_ _319_ _121_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__558__A1 _204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_602_ Datapath.k\[11\] Datapath.k\[10\] _248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__549__A1 _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_533_ _181_ _176_ _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_464_ _129_ _062_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_395_ _067_ _068_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_516_ _097_ _168_ _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_447_ _115_ Datapath.i\[4\] _062_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_378_ net18 _056_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__498__B _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__391__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__373__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__716__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I co[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__739__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__594__A2 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_695_ _329_ _333_ _334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I co[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_480_ _131_ _053_ _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__567__A2 _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_678_ _047_ Datapath.k\[16\] Datapath.k\[17\] _060_ _319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__558__A2 _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_601_ _246_ _247_ _080_ _158_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__549__A2 _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_532_ _182_ _183_ _184_ _158_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_394_ net12 net13 net14 net15 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_463_ _128_ Datapath.i\[7\] _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__485__A1 _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__467__A1 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_515_ _167_ _097_ _168_ _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_377_ Datapath.i\[12\] _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_446_ _113_ _114_ _115_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__689__B Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__612__A1 _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_429_ _102_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__603__A1 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 co[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__530__B1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__348__I _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__512__B1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_694_ _332_ _333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_677_ _313_ _315_ _317_ _318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__729__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_531_ Datapath.k\[4\] _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_600_ Datapath.k\[11\] _103_ _038_ net2 _046_ _247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_393_ net16 net2 net3 net4 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_462_ _126_ _128_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__485__A2 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_729_ _022_ clknet_2_2__leaf_clk Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__400__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__467__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_514_ Datapath.k\[3\] Datapath.k\[2\] _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_376_ net18 _055_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_445_ _113_ _045_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__458__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__612__A2 _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__376__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_428_ _073_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_359_ _041_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 co[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__358__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__530__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__588__A1 _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__512__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_693_ _330_ _331_ _332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__503__A1 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_676_ _316_ _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__552__I Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__494__A3 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_530_ net11 _120_ Datapath.k\[5\] _102_ _042_ _183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_461_ _127_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_392_ net1 _062_ _063_ _066_ FSM.NS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_728_ _021_ clknet_2_2__leaf_clk Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_659_ _284_ _293_ _300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_444_ _062_ Datapath.i\[3\] _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_513_ _165_ _162_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__719__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_375_ Datapath.i\[11\] _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__I Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_358_ net18 _045_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__376__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_427_ _065_ _094_ _097_ _100_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 co[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__530__A2 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__588__A2 _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_692_ Datapath.k\[18\] Datapath.k\[17\] _331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__503__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__375__I Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input14_I co[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_744_ FSM.NS\[1\] clknet_2_1__leaf_clk FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_675_ _036_ _037_ _316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__488__A1 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I co[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__651__A1 _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__403__A1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_460_ _125_ Datapath.i\[6\] _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_391_ _064_ _065_ _037_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_727_ _020_ clknet_2_2__leaf_clk Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_589_ Datapath.k\[10\] _103_ _038_ net16 _046_ _237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_658_ _297_ _298_ _299_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__633__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__563__I Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__624__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_512_ _160_ _166_ _096_ _158_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_443_ _110_ _037_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_374_ _054_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__551__B1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_357_ Datapath.i\[3\] _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_426_ _098_ _099_ _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput4 co[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__709__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_409_ Datapath.k\[16\] _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__504__C _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_691_ Datapath.k\[18\] Datapath.k\[17\] _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__430__B _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_743_ FSM.NS\[0\] clknet_2_3__leaf_clk FSM.CS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_674_ _304_ _308_ _314_ _315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__476__I _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__479__A2 _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__403__A2 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_390_ Datapath.k\[1\] _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_726_ _019_ clknet_2_2__leaf_clk Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_657_ _039_ Datapath.k\[15\] _299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_588_ _231_ _234_ _235_ _236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__397__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__742__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_511_ _164_ _036_ _165_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_442_ _112_ _044_ _109_ _106_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_373_ _047_ Datapath.i\[10\] _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__388__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__560__A1 _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_709_ _002_ clknet_2_0__leaf_clk Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__551__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__533__A1 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_356_ _044_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_425_ Datapath.k\[12\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 co[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_32_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__569__I _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_408_ Datapath.k\[17\] _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__506__A1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__389__I _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_690_ _309_ _327_ _328_ _329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__497__A3 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_742_ _035_ clknet_2_3__leaf_clk Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_673_ _312_ _314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_587_ _231_ _234_ _060_ _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_725_ _018_ clknet_2_2__leaf_clk Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_656_ Datapath.k\[16\] _103_ _038_ net7 _042_ _298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__609__B1 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_441_ _111_ _037_ _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_510_ _161_ Datapath.k\[0\] _162_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__388__A2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_372_ net18 _053_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__560__A2 _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_708_ _001_ clknet_2_0__leaf_clk Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_639_ _089_ _098_ _282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__551__A2 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_424_ Datapath.k\[13\] _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__533__A2 _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_355_ _042_ Datapath.i\[2\] _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__732__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 co[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__608__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__515__A2 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_407_ _079_ _080_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__506__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__681__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__433__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_741_ _034_ clknet_2_3__leaf_clk Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_672_ _309_ _312_ _313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__590__B1 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__581__B1 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I co[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_724_ _017_ clknet_2_1__leaf_clk Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_586_ _233_ _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_655_ _295_ _296_ _064_ _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__618__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I co[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__609__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__537__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_440_ _110_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_371_ Datapath.i\[9\] _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__560__A3 _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_707_ _000_ clknet_2_0__leaf_clk Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_569_ _215_ _218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__447__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_638_ _278_ _280_ _281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_423_ _095_ _096_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_354_ _043_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 co[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__515__A3 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__A2 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_406_ Datapath.k\[10\] _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__681__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__433__A2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__722__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 co[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_740_ _033_ clknet_2_3__leaf_clk Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_671_ _310_ _311_ _312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__590__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__645__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__581__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__632__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__572__A1 _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__627__A2 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_723_ _016_ clknet_2_3__leaf_clk Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_654_ _286_ _283_ _293_ _296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_585_ _077_ _232_ _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__618__A2 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__554__A1 _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_370_ net18 _052_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_637_ _279_ _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_706_ _341_ _342_ _343_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_568_ _175_ _216_ _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_499_ _064_ net1 _155_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__527__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_353_ _042_ Datapath.i\[1\] _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_422_ Datapath.k\[2\] _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_5_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 co[1] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_405_ Datapath.k\[11\] _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 co[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_670_ Datapath.k\[16\] Datapath.k\[15\] _311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__581__A2 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__712__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__572__A2 _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_653_ _290_ _291_ _294_ _295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_722_ _015_ clknet_2_0__leaf_clk Datapath.i\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_584_ Datapath.k\[9\] Datapath.k\[8\] _232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__735__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__554__A2 _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__481__A1 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_567_ _214_ _215_ _216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_636_ _263_ _271_ _279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_705_ _047_ Datapath.k\[19\] _343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_498_ _060_ Datapath.k\[0\] _037_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__527__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_421_ Datapath.k\[3\] _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__463__A1 _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_352_ _041_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 co[2] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__454__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_619_ _261_ _262_ _263_ _264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_404_ Datapath.k\[19\] Datapath.k\[18\] _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__675__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__427__A1 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__469__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__657__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 co[5] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__646__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__501__I _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_652_ _293_ _294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_721_ _014_ clknet_2_1__leaf_clk Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_583_ _227_ _224_ _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__539__B1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I co[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__490__A2 _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_704_ _335_ _331_ _339_ _342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__481__A2 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_566_ _198_ _207_ _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_635_ _257_ _259_ _277_ _278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_497_ _153_ _154_ _121_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_8_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I co[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__463__A2 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_420_ _093_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_351_ _039_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__725__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__454__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_549_ _194_ _198_ _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_618_ Datapath.k\[12\] Datapath.k\[11\] _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_403_ _075_ _076_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__372__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__675__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__427__A2 _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__363__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__414__I Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__657__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 co[6] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__584__A1 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__575__A1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__409__I Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__566__A1 _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__557__A1 _206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_720_ _013_ clknet_2_2__leaf_clk Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__548__A1 _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_582_ _229_ _230_ _076_ _158_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_651_ _090_ _292_ _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__539__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__422__I Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_703_ _340_ _317_ _341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_634_ _265_ _272_ _277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__481__A3 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_496_ _149_ _059_ _058_ _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_565_ _188_ _179_ _214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__417__I _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_350_ net18 _040_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_617_ _099_ _079_ _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_479_ _134_ _138_ _141_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_548_ _194_ _198_ _199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__678__B1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_402_ Datapath.k\[8\] _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__372__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__427__A3 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__363__A2 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__715__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 co[7] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__738__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__584__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__575__A2 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__425__I Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__566__A2 _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__557__A2 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_650_ Datapath.k\[15\] Datapath.k\[14\] _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__548__A2 _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_581_ net15 _120_ Datapath.k\[9\] _102_ _046_ _230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__484__A1 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__539__A2 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__466__A1 _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_702_ _335_ _331_ _339_ _340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_633_ _275_ _276_ _098_ _047_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_564_ _211_ _212_ _213_ _158_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_495_ _152_ Datapath.i\[15\] _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__679__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_547_ _196_ _197_ _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_616_ _260_ _261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_478_ _140_ _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__678__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__678__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__602__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_401_ Datapath.k\[9\] _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__427__A4 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 co[8] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__531__I Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__687__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__351__I _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__728__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_580_ _227_ _064_ _228_ _229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__484__A2 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__346__I _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__475__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__466__A2 Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_563_ Datapath.k\[7\] _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_632_ Datapath.k\[14\] _103_ _038_ net5 _046_ _276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_701_ _078_ _338_ _339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_494_ _151_ _152_ _121_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_5_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__448__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__384__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__589__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_546_ Datapath.k\[6\] Datapath.k\[5\] _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_615_ _257_ _259_ _260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_477_ _139_ Datapath.i\[10\] _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__678__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__534__I Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__366__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_400_ _072_ _039_ _073_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_529_ _180_ _064_ _181_ _182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__520__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__587__A1 _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 co[9] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__502__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__349__I Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__452__I _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__705__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__632__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__466__A3 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_700_ Datapath.k\[19\] Datapath.k\[18\] _338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__623__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_562_ net14 _120_ Datapath.k\[8\] _102_ _046_ _212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_493_ _149_ _058_ _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_631_ _273_ _274_ _036_ _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__718__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_614_ _258_ _242_ _248_ _259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_476_ _138_ _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_545_ _195_ _196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_459_ _125_ Datapath.i\[6\] _062_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_528_ _175_ _179_ _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__587__A2 _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__545__I _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__511__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 st net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__487__A1 _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__411__A1 _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__650__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__469__A1 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__632__B2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_630_ _270_ _272_ _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__623__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_561_ _208_ _064_ _210_ _211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_492_ _149_ _058_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_613_ _255_ _239_ _258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_475_ _135_ _037_ _123_ _137_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_544_ Datapath.k\[6\] Datapath.k\[5\] _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__532__B1 _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_527_ _175_ _179_ _180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__708__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_458_ _119_ _121_ _125_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_389_ _036_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__505__B1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__511__A3 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__556__I _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__487__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__411__A2 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__469__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__396__A1 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__632__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__623__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_560_ _200_ _195_ _209_ _210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_491_ _150_ _121_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__741__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_689_ Datapath.k\[17\] Datapath.k\[15\] Datapath.k\[16\] _328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__378__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__393__A4 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__605__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__541__A1 _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_543_ _181_ _193_ _087_ _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_612_ _217_ _220_ _256_ _257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_474_ _136_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__532__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__523__A1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__514__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_526_ _177_ _178_ _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__505__B2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_457_ _113_ _124_ _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ _047_ net17 _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__600__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_509_ _163_ _086_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__505__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__B Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__411__A3 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I st vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input9_I co[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__387__I _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__396__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__608__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_490_ Datapath.i\[13\] _146_ _149_ _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__378__A2 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_688_ _314_ _084_ _321_ _327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__550__A2 _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_611_ _238_ _255_ _256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_542_ _192_ _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_473_ Datapath.i\[9\] Datapath.i\[8\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__599__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__523__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__731__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__514__A2 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_525_ Datapath.k\[4\] Datapath.k\[3\] _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_456_ _123_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_387_ _061_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__505__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__432__A1 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__499__A1 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_439_ _106_ _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_508_ _161_ _162_ _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__562__B1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__396__A3 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__553__B1 _203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__608__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__578__I _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_687_ _325_ _326_ _121_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__550__A3 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_610_ _243_ _249_ _255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_541_ _186_ _095_ _184_ _192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_472_ _111_ _051_ _050_ _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_739_ _032_ clknet_2_3__leaf_clk Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_524_ _176_ _177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_455_ _122_ _045_ _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_386_ _038_ _060_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__441__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__586__I _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__519__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__432__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__499__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__423__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_438_ Datapath.i\[2\] _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_369_ Datapath.i\[8\] _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_507_ Datapath.k\[2\] Datapath.k\[1\] _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__721__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__350__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__744__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__580__A1 _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__399__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__562__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__617__A2 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__396__A4 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__553__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__608__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__544__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_686_ _042_ Datapath.k\[17\] Datapath.k\[18\] _060_ _326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__535__A1 _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_540_ _190_ _191_ _186_ _158_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_471_ _062_ Datapath.i\[10\] _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__517__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_738_ _031_ clknet_2_3__leaf_clk Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_669_ _083_ _088_ _310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_523_ Datapath.k\[4\] Datapath.k\[3\] _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_454_ Datapath.i\[5\] Datapath.i\[4\] _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_385_ FSM.CS\[0\] _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_506_ _096_ _065_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_437_ _043_ _107_ _108_ _040_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_368_ net18 _051_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__350__A2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__580__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__399__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__711__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__562__A2 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__734__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I co[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__544__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__480__A1 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_685_ _322_ _317_ _324_ _325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__535__A2 _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input7_I co[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__471__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__526__A2 _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_470_ _053_ _131_ _133_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__517__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_737_ _030_ clknet_2_3__leaf_clk Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_599_ _244_ _064_ _245_ _246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_668_ _304_ _308_ _309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__508__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__444__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_453_ _120_ _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_522_ _165_ _170_ _174_ _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_384_ _039_ _059_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__674__A1 _304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__459__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__551__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__656__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__656__B2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_436_ Datapath.i\[1\] _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_505_ net9 _121_ Datapath.k\[3\] _103_ _042_ _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_367_ Datapath.i\[7\] _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__647__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_419_ Datapath.k\[7\] Datapath.k\[6\] _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__401__I Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__480__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_684_ _315_ _311_ _323_ _324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__471__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__462__A2 _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__517__A3 _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_736_ _029_ clknet_2_3__leaf_clk Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_598_ _240_ _243_ _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_667_ _305_ _307_ _308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__724__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__692__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__380__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__435__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_452_ _061_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_521_ Datapath.k\[3\] Datapath.k\[1\] Datapath.k\[2\] _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_383_ Datapath.i\[15\] _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__674__A2 _308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_719_ _012_ clknet_2_2__leaf_clk Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__353__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_435_ _106_ _037_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_366_ net18 _050_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_504_ _060_ _065_ _096_ _073_ _159_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__583__A1 _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__574__A1 _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__562__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__565__A1 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_349_ Datapath.i\[0\] _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _085_ _086_ _087_ _091_ _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__538__A1 _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__701__A1 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_683_ _084_ _321_ _323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_735_ _028_ clknet_2_3__leaf_clk Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_597_ _240_ _243_ _244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_666_ _300_ _279_ _306_ _307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_520_ _172_ _173_ _095_ _158_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_382_ _039_ _058_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_451_ _118_ Datapath.i\[5\] _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_649_ _283_ _291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_718_ _011_ clknet_2_0__leaf_clk Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__420__I _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__714__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_503_ _121_ net8 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_434_ Datapath.i\[1\] Datapath.i\[0\] _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_365_ Datapath.i\[6\] _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__737__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__574__A2 _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__565__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _039_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_417_ _090_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__483__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__538__A2 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__529__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__465__A1 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_682_ _320_ _084_ _321_ _322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I co[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__686__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__686__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_734_ _027_ clknet_2_2__leaf_clk Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_665_ _283_ _292_ _306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_596_ _241_ _242_ _243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I co[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__601__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__668__A1 _304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_450_ _116_ _118_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_381_ Datapath.i\[14\] _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__581__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_648_ _278_ _280_ _284_ _290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_717_ _010_ clknet_2_0__leaf_clk Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_579_ _222_ _225_ _228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_433_ _039_ _040_ _105_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_502_ _156_ _157_ _086_ _158_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_364_ _049_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__587__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_416_ _088_ _089_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_347_ _036_ _038_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_24_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__727__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__529__A3 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_681_ Datapath.k\[17\] Datapath.k\[16\] _321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__392__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__447__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__686__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_733_ _026_ clknet_2_2__leaf_clk Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_595_ Datapath.k\[10\] Datapath.k\[9\] _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_664_ _259_ _302_ _305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__524__I _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__668__A2 _308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ net18 _057_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 x[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_716_ _009_ clknet_2_0__leaf_clk Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_578_ _226_ _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_647_ _288_ _289_ _089_ _047_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__347__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

