magic
tech gf180mcuC
magscale 1 10
timestamp 1670118490
<< metal1 >>
rect 1344 40794 42560 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 42560 40794
rect 1344 40708 42560 40742
rect 1344 40010 42560 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 42560 40010
rect 1344 39924 42560 39958
rect 1344 39226 42560 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 42560 39226
rect 1344 39140 42560 39174
rect 1344 38442 42560 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 42560 38442
rect 1344 38356 42560 38390
rect 1344 37658 42560 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 42560 37658
rect 1344 37572 42560 37606
rect 1344 36874 42560 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 42560 36874
rect 1344 36788 42560 36822
rect 1344 36090 42560 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 42560 36090
rect 1344 36004 42560 36038
rect 1344 35306 42560 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 42560 35306
rect 1344 35220 42560 35254
rect 1344 34522 42560 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 42560 34522
rect 1344 34436 42560 34470
rect 1344 33738 42560 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 42560 33738
rect 1344 33652 42560 33686
rect 1344 32954 42560 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 42560 32954
rect 1344 32868 42560 32902
rect 1344 32170 42560 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 42560 32170
rect 1344 32084 42560 32118
rect 1344 31386 42560 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 42560 31386
rect 1344 31300 42560 31334
rect 1344 30602 42560 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 42560 30602
rect 1344 30516 42560 30550
rect 1344 29818 42560 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 42560 29818
rect 1344 29732 42560 29766
rect 1344 29034 42560 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 42560 29034
rect 1344 28948 42560 28982
rect 1344 28250 42560 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 42560 28250
rect 1344 28164 42560 28198
rect 1344 27466 42560 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 42560 27466
rect 1344 27380 42560 27414
rect 1344 26682 42560 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 42560 26682
rect 1344 26596 42560 26630
rect 1344 25898 42560 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 42560 25898
rect 1344 25812 42560 25846
rect 2494 25506 2546 25518
rect 2494 25442 2546 25454
rect 2942 25282 2994 25294
rect 2942 25218 2994 25230
rect 5070 25282 5122 25294
rect 5070 25218 5122 25230
rect 5742 25282 5794 25294
rect 5742 25218 5794 25230
rect 6190 25282 6242 25294
rect 6190 25218 6242 25230
rect 6974 25282 7026 25294
rect 6974 25218 7026 25230
rect 7422 25282 7474 25294
rect 7422 25218 7474 25230
rect 7870 25282 7922 25294
rect 7870 25218 7922 25230
rect 9550 25282 9602 25294
rect 9550 25218 9602 25230
rect 1344 25114 42560 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 42560 25114
rect 1344 25028 42560 25062
rect 2270 24722 2322 24734
rect 2270 24658 2322 24670
rect 6862 24722 6914 24734
rect 6862 24658 6914 24670
rect 1822 24610 1874 24622
rect 1822 24546 1874 24558
rect 2718 24610 2770 24622
rect 2718 24546 2770 24558
rect 3278 24610 3330 24622
rect 3278 24546 3330 24558
rect 4062 24610 4114 24622
rect 4062 24546 4114 24558
rect 4510 24610 4562 24622
rect 4510 24546 4562 24558
rect 5070 24610 5122 24622
rect 5070 24546 5122 24558
rect 5518 24610 5570 24622
rect 5518 24546 5570 24558
rect 5966 24610 6018 24622
rect 5966 24546 6018 24558
rect 6414 24610 6466 24622
rect 6414 24546 6466 24558
rect 7310 24610 7362 24622
rect 7310 24546 7362 24558
rect 7646 24610 7698 24622
rect 7646 24546 7698 24558
rect 8206 24610 8258 24622
rect 8206 24546 8258 24558
rect 8654 24610 8706 24622
rect 8654 24546 8706 24558
rect 9102 24610 9154 24622
rect 9102 24546 9154 24558
rect 9998 24610 10050 24622
rect 9998 24546 10050 24558
rect 10670 24610 10722 24622
rect 10670 24546 10722 24558
rect 11118 24610 11170 24622
rect 11118 24546 11170 24558
rect 8082 24446 8094 24498
rect 8146 24495 8158 24498
rect 9090 24495 9102 24498
rect 8146 24449 9102 24495
rect 8146 24446 8158 24449
rect 9090 24446 9102 24449
rect 9154 24446 9166 24498
rect 1344 24330 42560 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 42560 24330
rect 1344 24244 42560 24278
rect 8754 24110 8766 24162
rect 8818 24159 8830 24162
rect 9538 24159 9550 24162
rect 8818 24113 9550 24159
rect 8818 24110 8830 24113
rect 9538 24110 9550 24113
rect 9602 24110 9614 24162
rect 8654 24050 8706 24062
rect 8654 23986 8706 23998
rect 9102 24050 9154 24062
rect 9102 23986 9154 23998
rect 11230 24050 11282 24062
rect 11230 23986 11282 23998
rect 12238 24050 12290 24062
rect 12238 23986 12290 23998
rect 14030 24050 14082 24062
rect 14030 23986 14082 23998
rect 14478 24050 14530 24062
rect 14478 23986 14530 23998
rect 15038 24050 15090 24062
rect 15038 23986 15090 23998
rect 13582 23938 13634 23950
rect 13582 23874 13634 23886
rect 3726 23826 3778 23838
rect 3726 23762 3778 23774
rect 5742 23826 5794 23838
rect 5742 23762 5794 23774
rect 8318 23826 8370 23838
rect 8318 23762 8370 23774
rect 1934 23714 1986 23726
rect 1934 23650 1986 23662
rect 2382 23714 2434 23726
rect 2382 23650 2434 23662
rect 2830 23714 2882 23726
rect 2830 23650 2882 23662
rect 3278 23714 3330 23726
rect 3278 23650 3330 23662
rect 4174 23714 4226 23726
rect 4174 23650 4226 23662
rect 4622 23714 4674 23726
rect 4622 23650 4674 23662
rect 4958 23714 5010 23726
rect 4958 23650 5010 23662
rect 6302 23714 6354 23726
rect 6302 23650 6354 23662
rect 6862 23714 6914 23726
rect 6862 23650 6914 23662
rect 7422 23714 7474 23726
rect 7422 23650 7474 23662
rect 7758 23714 7810 23726
rect 7758 23650 7810 23662
rect 9662 23714 9714 23726
rect 9662 23650 9714 23662
rect 10110 23714 10162 23726
rect 10110 23650 10162 23662
rect 10894 23714 10946 23726
rect 10894 23650 10946 23662
rect 11902 23714 11954 23726
rect 11902 23650 11954 23662
rect 12686 23714 12738 23726
rect 12686 23650 12738 23662
rect 1344 23546 42560 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 42560 23546
rect 1344 23460 42560 23494
rect 2158 23378 2210 23390
rect 2158 23314 2210 23326
rect 10222 23154 10274 23166
rect 10222 23090 10274 23102
rect 13022 23154 13074 23166
rect 13022 23090 13074 23102
rect 16830 23154 16882 23166
rect 16830 23090 16882 23102
rect 1822 23042 1874 23054
rect 1822 22978 1874 22990
rect 2606 23042 2658 23054
rect 2606 22978 2658 22990
rect 3166 23042 3218 23054
rect 3166 22978 3218 22990
rect 3614 23042 3666 23054
rect 3614 22978 3666 22990
rect 3950 23042 4002 23054
rect 3950 22978 4002 22990
rect 4398 23042 4450 23054
rect 4398 22978 4450 22990
rect 4846 23042 4898 23054
rect 4846 22978 4898 22990
rect 5518 23042 5570 23054
rect 5518 22978 5570 22990
rect 6190 23042 6242 23054
rect 6190 22978 6242 22990
rect 6526 23042 6578 23054
rect 6526 22978 6578 22990
rect 7086 23042 7138 23054
rect 7086 22978 7138 22990
rect 7422 23042 7474 23054
rect 7422 22978 7474 22990
rect 7870 23042 7922 23054
rect 7870 22978 7922 22990
rect 8542 23042 8594 23054
rect 8542 22978 8594 22990
rect 9102 23042 9154 23054
rect 9102 22978 9154 22990
rect 9662 23042 9714 23054
rect 9662 22978 9714 22990
rect 10670 23042 10722 23054
rect 10670 22978 10722 22990
rect 11342 23042 11394 23054
rect 11342 22978 11394 22990
rect 12014 23042 12066 23054
rect 12014 22978 12066 22990
rect 12462 23042 12514 23054
rect 12462 22978 12514 22990
rect 13470 23042 13522 23054
rect 13470 22978 13522 22990
rect 13806 23042 13858 23054
rect 13806 22978 13858 22990
rect 14702 23042 14754 23054
rect 14702 22978 14754 22990
rect 15150 23042 15202 23054
rect 15150 22978 15202 22990
rect 15486 23042 15538 23054
rect 15486 22978 15538 22990
rect 16046 23042 16098 23054
rect 16046 22978 16098 22990
rect 16494 23042 16546 23054
rect 16494 22978 16546 22990
rect 1344 22762 42560 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 42560 22762
rect 1344 22676 42560 22710
rect 3938 22542 3950 22594
rect 4002 22591 4014 22594
rect 4946 22591 4958 22594
rect 4002 22545 4958 22591
rect 4002 22542 4014 22545
rect 4946 22542 4958 22545
rect 5010 22542 5022 22594
rect 1822 22482 1874 22494
rect 1822 22418 1874 22430
rect 2718 22482 2770 22494
rect 2718 22418 2770 22430
rect 3054 22482 3106 22494
rect 3054 22418 3106 22430
rect 4398 22482 4450 22494
rect 4398 22418 4450 22430
rect 4846 22482 4898 22494
rect 4846 22418 4898 22430
rect 11342 22482 11394 22494
rect 11342 22418 11394 22430
rect 17390 22482 17442 22494
rect 17390 22418 17442 22430
rect 17838 22482 17890 22494
rect 17838 22418 17890 22430
rect 39106 22318 39118 22370
rect 39170 22318 39182 22370
rect 10110 22258 10162 22270
rect 10110 22194 10162 22206
rect 16494 22258 16546 22270
rect 40002 22206 40014 22258
rect 40066 22206 40078 22258
rect 16494 22194 16546 22206
rect 2158 22146 2210 22158
rect 2158 22082 2210 22094
rect 3614 22146 3666 22158
rect 3614 22082 3666 22094
rect 4062 22146 4114 22158
rect 4062 22082 4114 22094
rect 6078 22146 6130 22158
rect 6078 22082 6130 22094
rect 6414 22146 6466 22158
rect 6414 22082 6466 22094
rect 6862 22146 6914 22158
rect 6862 22082 6914 22094
rect 7758 22146 7810 22158
rect 7758 22082 7810 22094
rect 8094 22146 8146 22158
rect 8094 22082 8146 22094
rect 8542 22146 8594 22158
rect 8542 22082 8594 22094
rect 8990 22146 9042 22158
rect 8990 22082 9042 22094
rect 9550 22146 9602 22158
rect 9550 22082 9602 22094
rect 10446 22146 10498 22158
rect 10446 22082 10498 22094
rect 11006 22146 11058 22158
rect 11006 22082 11058 22094
rect 11790 22146 11842 22158
rect 11790 22082 11842 22094
rect 12350 22146 12402 22158
rect 12350 22082 12402 22094
rect 12910 22146 12962 22158
rect 12910 22082 12962 22094
rect 13694 22146 13746 22158
rect 13694 22082 13746 22094
rect 14142 22146 14194 22158
rect 14142 22082 14194 22094
rect 14926 22146 14978 22158
rect 14926 22082 14978 22094
rect 15374 22146 15426 22158
rect 15374 22082 15426 22094
rect 16158 22146 16210 22158
rect 16158 22082 16210 22094
rect 16942 22146 16994 22158
rect 16942 22082 16994 22094
rect 18286 22146 18338 22158
rect 18286 22082 18338 22094
rect 40574 22146 40626 22158
rect 40574 22082 40626 22094
rect 1344 21978 42560 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 42560 21978
rect 1344 21892 42560 21926
rect 2942 21810 2994 21822
rect 2942 21746 2994 21758
rect 4734 21810 4786 21822
rect 4734 21746 4786 21758
rect 5742 21810 5794 21822
rect 5742 21746 5794 21758
rect 6190 21810 6242 21822
rect 6190 21746 6242 21758
rect 7982 21810 8034 21822
rect 7982 21746 8034 21758
rect 10110 21810 10162 21822
rect 10110 21746 10162 21758
rect 10558 21810 10610 21822
rect 10558 21746 10610 21758
rect 11006 21810 11058 21822
rect 11006 21746 11058 21758
rect 14030 21810 14082 21822
rect 14030 21746 14082 21758
rect 16942 21810 16994 21822
rect 16942 21746 16994 21758
rect 17614 21810 17666 21822
rect 17614 21746 17666 21758
rect 19406 21810 19458 21822
rect 19406 21746 19458 21758
rect 4286 21698 4338 21710
rect 4286 21634 4338 21646
rect 16046 21698 16098 21710
rect 16046 21634 16098 21646
rect 16494 21698 16546 21710
rect 16494 21634 16546 21646
rect 3838 21586 3890 21598
rect 3838 21522 3890 21534
rect 5406 21586 5458 21598
rect 5406 21522 5458 21534
rect 2158 21474 2210 21486
rect 2158 21410 2210 21422
rect 2606 21474 2658 21486
rect 2606 21410 2658 21422
rect 3502 21474 3554 21486
rect 3502 21410 3554 21422
rect 6750 21474 6802 21486
rect 6750 21410 6802 21422
rect 7086 21474 7138 21486
rect 7086 21410 7138 21422
rect 7534 21474 7586 21486
rect 7534 21410 7586 21422
rect 8542 21474 8594 21486
rect 8542 21410 8594 21422
rect 9102 21474 9154 21486
rect 9102 21410 9154 21422
rect 9662 21474 9714 21486
rect 9662 21410 9714 21422
rect 11454 21474 11506 21486
rect 11454 21410 11506 21422
rect 12014 21474 12066 21486
rect 12014 21410 12066 21422
rect 12350 21474 12402 21486
rect 12350 21410 12402 21422
rect 13246 21474 13298 21486
rect 13246 21410 13298 21422
rect 13694 21474 13746 21486
rect 13694 21410 13746 21422
rect 14478 21474 14530 21486
rect 14478 21410 14530 21422
rect 14926 21474 14978 21486
rect 14926 21410 14978 21422
rect 15598 21474 15650 21486
rect 15598 21410 15650 21422
rect 18174 21474 18226 21486
rect 18174 21410 18226 21422
rect 18510 21474 18562 21486
rect 18510 21410 18562 21422
rect 18958 21474 19010 21486
rect 18958 21410 19010 21422
rect 2818 21310 2830 21362
rect 2882 21359 2894 21362
rect 3602 21359 3614 21362
rect 2882 21313 3614 21359
rect 2882 21310 2894 21313
rect 3602 21310 3614 21313
rect 3666 21310 3678 21362
rect 8530 21310 8542 21362
rect 8594 21359 8606 21362
rect 8866 21359 8878 21362
rect 8594 21313 8878 21359
rect 8594 21310 8606 21313
rect 8866 21310 8878 21313
rect 8930 21310 8942 21362
rect 9650 21310 9662 21362
rect 9714 21359 9726 21362
rect 10770 21359 10782 21362
rect 9714 21313 10782 21359
rect 9714 21310 9726 21313
rect 10770 21310 10782 21313
rect 10834 21359 10846 21362
rect 11442 21359 11454 21362
rect 10834 21313 11454 21359
rect 10834 21310 10846 21313
rect 11442 21310 11454 21313
rect 11506 21359 11518 21362
rect 12338 21359 12350 21362
rect 11506 21313 12350 21359
rect 11506 21310 11518 21313
rect 12338 21310 12350 21313
rect 12402 21310 12414 21362
rect 1344 21194 42560 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 42560 21194
rect 1344 21108 42560 21142
rect 1922 20974 1934 21026
rect 1986 21023 1998 21026
rect 2482 21023 2494 21026
rect 1986 20977 2494 21023
rect 1986 20974 1998 20977
rect 2482 20974 2494 20977
rect 2546 20974 2558 21026
rect 13794 20974 13806 21026
rect 13858 21023 13870 21026
rect 14578 21023 14590 21026
rect 13858 20977 14590 21023
rect 13858 20974 13870 20977
rect 14578 20974 14590 20977
rect 14642 20974 14654 21026
rect 2382 20914 2434 20926
rect 2382 20850 2434 20862
rect 5630 20914 5682 20926
rect 5630 20850 5682 20862
rect 7086 20914 7138 20926
rect 7086 20850 7138 20862
rect 8990 20914 9042 20926
rect 8990 20850 9042 20862
rect 11902 20914 11954 20926
rect 11902 20850 11954 20862
rect 2046 20690 2098 20702
rect 2046 20626 2098 20638
rect 7982 20690 8034 20702
rect 7982 20626 8034 20638
rect 19630 20690 19682 20702
rect 19630 20626 19682 20638
rect 2830 20578 2882 20590
rect 2830 20514 2882 20526
rect 3502 20578 3554 20590
rect 3502 20514 3554 20526
rect 3950 20578 4002 20590
rect 3950 20514 4002 20526
rect 4622 20578 4674 20590
rect 4622 20514 4674 20526
rect 5070 20578 5122 20590
rect 5070 20514 5122 20526
rect 6302 20578 6354 20590
rect 6302 20514 6354 20526
rect 6638 20578 6690 20590
rect 6638 20514 6690 20526
rect 7646 20578 7698 20590
rect 7646 20514 7698 20526
rect 8542 20578 8594 20590
rect 8542 20514 8594 20526
rect 9438 20578 9490 20590
rect 9438 20514 9490 20526
rect 10222 20578 10274 20590
rect 10222 20514 10274 20526
rect 10670 20578 10722 20590
rect 10670 20514 10722 20526
rect 11454 20578 11506 20590
rect 11454 20514 11506 20526
rect 12462 20578 12514 20590
rect 12462 20514 12514 20526
rect 12910 20578 12962 20590
rect 12910 20514 12962 20526
rect 13582 20578 13634 20590
rect 13582 20514 13634 20526
rect 14142 20578 14194 20590
rect 14142 20514 14194 20526
rect 14590 20578 14642 20590
rect 14590 20514 14642 20526
rect 15038 20578 15090 20590
rect 15038 20514 15090 20526
rect 15822 20578 15874 20590
rect 15822 20514 15874 20526
rect 16270 20578 16322 20590
rect 16270 20514 16322 20526
rect 16606 20578 16658 20590
rect 16606 20514 16658 20526
rect 17390 20578 17442 20590
rect 17390 20514 17442 20526
rect 17950 20578 18002 20590
rect 17950 20514 18002 20526
rect 18286 20578 18338 20590
rect 18286 20514 18338 20526
rect 18734 20578 18786 20590
rect 18734 20514 18786 20526
rect 19182 20578 19234 20590
rect 19182 20514 19234 20526
rect 20078 20578 20130 20590
rect 20078 20514 20130 20526
rect 1344 20410 42560 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 42560 20410
rect 1344 20324 42560 20358
rect 1934 20242 1986 20254
rect 1934 20178 1986 20190
rect 2718 20242 2770 20254
rect 2718 20178 2770 20190
rect 4734 20242 4786 20254
rect 4734 20178 4786 20190
rect 11342 20242 11394 20254
rect 11342 20178 11394 20190
rect 18286 20242 18338 20254
rect 18286 20178 18338 20190
rect 20526 20242 20578 20254
rect 20526 20178 20578 20190
rect 3166 20130 3218 20142
rect 3166 20066 3218 20078
rect 6750 20130 6802 20142
rect 6750 20066 6802 20078
rect 10894 20130 10946 20142
rect 10894 20066 10946 20078
rect 12462 20130 12514 20142
rect 12462 20066 12514 20078
rect 13358 20130 13410 20142
rect 13358 20066 13410 20078
rect 15038 20130 15090 20142
rect 15038 20066 15090 20078
rect 20974 20130 21026 20142
rect 20974 20066 21026 20078
rect 8542 20018 8594 20030
rect 8542 19954 8594 19966
rect 10446 20018 10498 20030
rect 10446 19954 10498 19966
rect 2270 19906 2322 19918
rect 2270 19842 2322 19854
rect 4062 19906 4114 19918
rect 4062 19842 4114 19854
rect 5182 19906 5234 19918
rect 5182 19842 5234 19854
rect 5966 19906 6018 19918
rect 5966 19842 6018 19854
rect 7198 19906 7250 19918
rect 7198 19842 7250 19854
rect 7646 19906 7698 19918
rect 7646 19842 7698 19854
rect 8206 19906 8258 19918
rect 8206 19842 8258 19854
rect 8990 19906 9042 19918
rect 8990 19842 9042 19854
rect 9662 19906 9714 19918
rect 9662 19842 9714 19854
rect 12014 19906 12066 19918
rect 12014 19842 12066 19854
rect 13022 19906 13074 19918
rect 13022 19842 13074 19854
rect 14030 19906 14082 19918
rect 14030 19842 14082 19854
rect 14478 19906 14530 19918
rect 14478 19842 14530 19854
rect 15598 19906 15650 19918
rect 15598 19842 15650 19854
rect 16046 19906 16098 19918
rect 16046 19842 16098 19854
rect 16718 19906 16770 19918
rect 16718 19842 16770 19854
rect 17950 19906 18002 19918
rect 17950 19842 18002 19854
rect 18734 19906 18786 19918
rect 18734 19842 18786 19854
rect 19294 19906 19346 19918
rect 19294 19842 19346 19854
rect 19630 19906 19682 19918
rect 19630 19842 19682 19854
rect 20078 19906 20130 19918
rect 20078 19842 20130 19854
rect 21422 19906 21474 19918
rect 21422 19842 21474 19854
rect 1698 19742 1710 19794
rect 1762 19791 1774 19794
rect 2258 19791 2270 19794
rect 1762 19745 2270 19791
rect 1762 19742 1774 19745
rect 2258 19742 2270 19745
rect 2322 19742 2334 19794
rect 7634 19742 7646 19794
rect 7698 19791 7710 19794
rect 8306 19791 8318 19794
rect 7698 19745 8318 19791
rect 7698 19742 7710 19745
rect 8306 19742 8318 19745
rect 8370 19742 8382 19794
rect 1344 19626 42560 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 42560 19626
rect 1344 19540 42560 19574
rect 9886 19458 9938 19470
rect 1810 19406 1822 19458
rect 1874 19455 1886 19458
rect 2818 19455 2830 19458
rect 1874 19409 2830 19455
rect 1874 19406 1886 19409
rect 2818 19406 2830 19409
rect 2882 19455 2894 19458
rect 3154 19455 3166 19458
rect 2882 19409 3166 19455
rect 2882 19406 2894 19409
rect 3154 19406 3166 19409
rect 3218 19406 3230 19458
rect 5730 19406 5742 19458
rect 5794 19455 5806 19458
rect 6178 19455 6190 19458
rect 5794 19409 6190 19455
rect 5794 19406 5806 19409
rect 6178 19406 6190 19409
rect 6242 19406 6254 19458
rect 7298 19406 7310 19458
rect 7362 19455 7374 19458
rect 7634 19455 7646 19458
rect 7362 19409 7646 19455
rect 7362 19406 7374 19409
rect 7634 19406 7646 19409
rect 7698 19406 7710 19458
rect 11330 19406 11342 19458
rect 11394 19455 11406 19458
rect 11554 19455 11566 19458
rect 11394 19409 11566 19455
rect 11394 19406 11406 19409
rect 11554 19406 11566 19409
rect 11618 19406 11630 19458
rect 12226 19406 12238 19458
rect 12290 19455 12302 19458
rect 12786 19455 12798 19458
rect 12290 19409 12798 19455
rect 12290 19406 12302 19409
rect 12786 19406 12798 19409
rect 12850 19406 12862 19458
rect 9886 19394 9938 19406
rect 1934 19346 1986 19358
rect 1934 19282 1986 19294
rect 3166 19346 3218 19358
rect 3166 19282 3218 19294
rect 4062 19346 4114 19358
rect 4062 19282 4114 19294
rect 5742 19346 5794 19358
rect 5742 19282 5794 19294
rect 7086 19346 7138 19358
rect 7086 19282 7138 19294
rect 13582 19346 13634 19358
rect 13582 19282 13634 19294
rect 18062 19346 18114 19358
rect 18062 19282 18114 19294
rect 19406 19346 19458 19358
rect 19406 19282 19458 19294
rect 20302 19346 20354 19358
rect 20302 19282 20354 19294
rect 22430 19346 22482 19358
rect 22430 19282 22482 19294
rect 9774 19234 9826 19246
rect 9774 19170 9826 19182
rect 10446 19234 10498 19246
rect 10446 19170 10498 19182
rect 11678 19234 11730 19246
rect 11678 19170 11730 19182
rect 2270 19122 2322 19134
rect 2270 19058 2322 19070
rect 7646 19122 7698 19134
rect 7646 19058 7698 19070
rect 8094 19122 8146 19134
rect 8094 19058 8146 19070
rect 8990 19122 9042 19134
rect 8990 19058 9042 19070
rect 9886 19122 9938 19134
rect 9886 19058 9938 19070
rect 18510 19122 18562 19134
rect 18510 19058 18562 19070
rect 18958 19122 19010 19134
rect 18958 19058 19010 19070
rect 2718 19010 2770 19022
rect 2718 18946 2770 18958
rect 3614 19010 3666 19022
rect 3614 18946 3666 18958
rect 4622 19010 4674 19022
rect 4622 18946 4674 18958
rect 5070 19010 5122 19022
rect 5070 18946 5122 18958
rect 6302 19010 6354 19022
rect 6302 18946 6354 18958
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 8206 19010 8258 19022
rect 8206 18946 8258 18958
rect 8878 19010 8930 19022
rect 8878 18946 8930 18958
rect 11230 19010 11282 19022
rect 11230 18946 11282 18958
rect 12238 19010 12290 19022
rect 12238 18946 12290 18958
rect 12686 19010 12738 19022
rect 12686 18946 12738 18958
rect 14142 19010 14194 19022
rect 14142 18946 14194 18958
rect 14702 19010 14754 19022
rect 14702 18946 14754 18958
rect 15150 19010 15202 19022
rect 15150 18946 15202 18958
rect 15598 19010 15650 19022
rect 15598 18946 15650 18958
rect 15934 19010 15986 19022
rect 15934 18946 15986 18958
rect 16606 19010 16658 19022
rect 16606 18946 16658 18958
rect 16942 19010 16994 19022
rect 16942 18946 16994 18958
rect 17390 19010 17442 19022
rect 17390 18946 17442 18958
rect 19854 19010 19906 19022
rect 19854 18946 19906 18958
rect 20750 19010 20802 19022
rect 20750 18946 20802 18958
rect 21534 19010 21586 19022
rect 21534 18946 21586 18958
rect 21982 19010 22034 19022
rect 21982 18946 22034 18958
rect 1344 18842 42560 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 42560 18842
rect 1344 18756 42560 18790
rect 3502 18674 3554 18686
rect 3502 18610 3554 18622
rect 4846 18674 4898 18686
rect 4846 18610 4898 18622
rect 7310 18674 7362 18686
rect 8878 18674 8930 18686
rect 7310 18610 7362 18622
rect 8094 18618 8146 18630
rect 6302 18562 6354 18574
rect 6302 18498 6354 18510
rect 6414 18562 6466 18574
rect 6414 18498 6466 18510
rect 7198 18562 7250 18574
rect 8878 18610 8930 18622
rect 9886 18674 9938 18686
rect 9886 18610 9938 18622
rect 10894 18674 10946 18686
rect 10894 18610 10946 18622
rect 11790 18674 11842 18686
rect 11790 18610 11842 18622
rect 12126 18674 12178 18686
rect 12126 18610 12178 18622
rect 12798 18674 12850 18686
rect 12798 18610 12850 18622
rect 22430 18674 22482 18686
rect 22430 18610 22482 18622
rect 8094 18554 8146 18566
rect 9774 18562 9826 18574
rect 7198 18498 7250 18510
rect 9774 18498 9826 18510
rect 11006 18562 11058 18574
rect 11006 18498 11058 18510
rect 12686 18562 12738 18574
rect 12686 18498 12738 18510
rect 1822 18450 1874 18462
rect 1822 18386 1874 18398
rect 6638 18450 6690 18462
rect 6638 18386 6690 18398
rect 7534 18450 7586 18462
rect 7534 18386 7586 18398
rect 7982 18450 8034 18462
rect 7982 18386 8034 18398
rect 8654 18450 8706 18462
rect 8654 18386 8706 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 14702 18450 14754 18462
rect 14702 18386 14754 18398
rect 17614 18450 17666 18462
rect 17614 18386 17666 18398
rect 18174 18450 18226 18462
rect 18174 18386 18226 18398
rect 19630 18450 19682 18462
rect 19630 18386 19682 18398
rect 22878 18450 22930 18462
rect 22878 18386 22930 18398
rect 2158 18338 2210 18350
rect 2158 18274 2210 18286
rect 2718 18338 2770 18350
rect 2718 18274 2770 18286
rect 3166 18338 3218 18350
rect 3166 18274 3218 18286
rect 3950 18338 4002 18350
rect 3950 18274 4002 18286
rect 4398 18338 4450 18350
rect 4398 18274 4450 18286
rect 5294 18338 5346 18350
rect 5294 18274 5346 18286
rect 5854 18338 5906 18350
rect 5854 18274 5906 18286
rect 13582 18338 13634 18350
rect 13582 18274 13634 18286
rect 14142 18338 14194 18350
rect 14142 18274 14194 18286
rect 15150 18338 15202 18350
rect 15150 18274 15202 18286
rect 15598 18338 15650 18350
rect 15598 18274 15650 18286
rect 16158 18338 16210 18350
rect 16158 18274 16210 18286
rect 16606 18338 16658 18350
rect 16606 18274 16658 18286
rect 18622 18338 18674 18350
rect 18622 18274 18674 18286
rect 19182 18338 19234 18350
rect 19182 18274 19234 18286
rect 20190 18338 20242 18350
rect 20190 18274 20242 18286
rect 20638 18338 20690 18350
rect 20638 18274 20690 18286
rect 21086 18338 21138 18350
rect 21086 18274 21138 18286
rect 21646 18338 21698 18350
rect 21646 18274 21698 18286
rect 21982 18338 22034 18350
rect 21982 18274 22034 18286
rect 8094 18226 8146 18238
rect 3602 18174 3614 18226
rect 3666 18223 3678 18226
rect 4386 18223 4398 18226
rect 3666 18177 4398 18223
rect 3666 18174 3678 18177
rect 4386 18174 4398 18177
rect 4450 18223 4462 18226
rect 6066 18223 6078 18226
rect 4450 18177 6078 18223
rect 4450 18174 4462 18177
rect 6066 18174 6078 18177
rect 6130 18174 6142 18226
rect 8094 18162 8146 18174
rect 9886 18226 9938 18238
rect 9886 18162 9938 18174
rect 10894 18226 10946 18238
rect 10894 18162 10946 18174
rect 12798 18226 12850 18238
rect 12798 18162 12850 18174
rect 13470 18226 13522 18238
rect 13470 18162 13522 18174
rect 14254 18226 14306 18238
rect 14578 18174 14590 18226
rect 14642 18223 14654 18226
rect 15026 18223 15038 18226
rect 14642 18177 15038 18223
rect 14642 18174 14654 18177
rect 15026 18174 15038 18177
rect 15090 18174 15102 18226
rect 15474 18174 15486 18226
rect 15538 18223 15550 18226
rect 16594 18223 16606 18226
rect 15538 18177 16606 18223
rect 15538 18174 15550 18177
rect 16594 18174 16606 18177
rect 16658 18174 16670 18226
rect 14254 18162 14306 18174
rect 1344 18058 42560 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 42560 18058
rect 1344 17972 42560 18006
rect 4062 17890 4114 17902
rect 4062 17826 4114 17838
rect 4846 17890 4898 17902
rect 4846 17826 4898 17838
rect 6302 17890 6354 17902
rect 6302 17826 6354 17838
rect 8430 17890 8482 17902
rect 18946 17838 18958 17890
rect 19010 17887 19022 17890
rect 19618 17887 19630 17890
rect 19010 17841 19630 17887
rect 19010 17838 19022 17841
rect 19618 17838 19630 17841
rect 19682 17838 19694 17890
rect 8430 17826 8482 17838
rect 2046 17778 2098 17790
rect 2046 17714 2098 17726
rect 3390 17778 3442 17790
rect 16830 17778 16882 17790
rect 9090 17726 9102 17778
rect 9154 17726 9166 17778
rect 3390 17714 3442 17726
rect 16830 17714 16882 17726
rect 17390 17778 17442 17790
rect 17390 17714 17442 17726
rect 18062 17778 18114 17790
rect 18062 17714 18114 17726
rect 18958 17778 19010 17790
rect 18958 17714 19010 17726
rect 22542 17778 22594 17790
rect 22542 17714 22594 17726
rect 23550 17778 23602 17790
rect 23550 17714 23602 17726
rect 2606 17666 2658 17678
rect 2606 17602 2658 17614
rect 5630 17666 5682 17678
rect 5630 17602 5682 17614
rect 6190 17666 6242 17678
rect 6190 17602 6242 17614
rect 7198 17666 7250 17678
rect 7198 17602 7250 17614
rect 7534 17666 7586 17678
rect 14702 17666 14754 17678
rect 12002 17614 12014 17666
rect 12066 17614 12078 17666
rect 12674 17614 12686 17666
rect 12738 17614 12750 17666
rect 7534 17602 7586 17614
rect 14702 17602 14754 17614
rect 15374 17666 15426 17678
rect 15374 17602 15426 17614
rect 3950 17554 4002 17566
rect 3950 17490 4002 17502
rect 4958 17554 5010 17566
rect 4958 17490 5010 17502
rect 6302 17554 6354 17566
rect 6302 17490 6354 17502
rect 8542 17554 8594 17566
rect 14030 17554 14082 17566
rect 11218 17502 11230 17554
rect 11282 17502 11294 17554
rect 8542 17490 8594 17502
rect 14030 17490 14082 17502
rect 14142 17554 14194 17566
rect 14142 17490 14194 17502
rect 3054 17442 3106 17454
rect 3054 17378 3106 17390
rect 4846 17442 4898 17454
rect 4846 17378 4898 17390
rect 7422 17442 7474 17454
rect 7422 17378 7474 17390
rect 8430 17442 8482 17454
rect 8430 17378 8482 17390
rect 12686 17442 12738 17454
rect 12686 17378 12738 17390
rect 13806 17442 13858 17454
rect 13806 17378 13858 17390
rect 14814 17442 14866 17454
rect 14814 17378 14866 17390
rect 15038 17442 15090 17454
rect 15038 17378 15090 17390
rect 16046 17442 16098 17454
rect 16046 17378 16098 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 19966 17442 20018 17454
rect 19966 17378 20018 17390
rect 20414 17442 20466 17454
rect 20414 17378 20466 17390
rect 20862 17442 20914 17454
rect 20862 17378 20914 17390
rect 21534 17442 21586 17454
rect 21534 17378 21586 17390
rect 22094 17442 22146 17454
rect 22094 17378 22146 17390
rect 23102 17442 23154 17454
rect 23102 17378 23154 17390
rect 24334 17442 24386 17454
rect 24334 17378 24386 17390
rect 26910 17442 26962 17454
rect 26910 17378 26962 17390
rect 1344 17274 42560 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 42560 17274
rect 1344 17188 42560 17222
rect 2046 17106 2098 17118
rect 2046 17042 2098 17054
rect 2830 17106 2882 17118
rect 2830 17042 2882 17054
rect 3054 17106 3106 17118
rect 3054 17042 3106 17054
rect 4510 17106 4562 17118
rect 4510 17042 4562 17054
rect 5294 17106 5346 17118
rect 5294 17042 5346 17054
rect 6190 17106 6242 17118
rect 6190 17042 6242 17054
rect 6974 17106 7026 17118
rect 6974 17042 7026 17054
rect 8430 17106 8482 17118
rect 8430 17042 8482 17054
rect 9102 17106 9154 17118
rect 9102 17042 9154 17054
rect 9662 17106 9714 17118
rect 9662 17042 9714 17054
rect 10334 17106 10386 17118
rect 10334 17042 10386 17054
rect 11566 17106 11618 17118
rect 11566 17042 11618 17054
rect 11678 17106 11730 17118
rect 11678 17042 11730 17054
rect 13582 17106 13634 17118
rect 13582 17042 13634 17054
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 19854 17106 19906 17118
rect 19854 17042 19906 17054
rect 22654 17106 22706 17118
rect 22654 17042 22706 17054
rect 23550 17106 23602 17118
rect 23550 17042 23602 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 1934 16994 1986 17006
rect 1934 16930 1986 16942
rect 2718 16994 2770 17006
rect 2718 16930 2770 16942
rect 3726 16994 3778 17006
rect 3726 16930 3778 16942
rect 4398 16994 4450 17006
rect 4398 16930 4450 16942
rect 5070 16994 5122 17006
rect 5070 16930 5122 16942
rect 5406 16994 5458 17006
rect 5406 16930 5458 16942
rect 6414 16994 6466 17006
rect 6414 16930 6466 16942
rect 6526 16994 6578 17006
rect 6526 16930 6578 16942
rect 7646 16994 7698 17006
rect 7646 16930 7698 16942
rect 8542 16994 8594 17006
rect 8542 16930 8594 16942
rect 10222 16994 10274 17006
rect 10222 16930 10274 16942
rect 11342 16994 11394 17006
rect 11342 16930 11394 16942
rect 11902 16994 11954 17006
rect 11902 16930 11954 16942
rect 12574 16994 12626 17006
rect 12574 16930 12626 16942
rect 12686 16994 12738 17006
rect 12686 16930 12738 16942
rect 13806 16994 13858 17006
rect 13806 16930 13858 16942
rect 17726 16994 17778 17006
rect 17726 16930 17778 16942
rect 18398 16994 18450 17006
rect 18398 16930 18450 16942
rect 18510 16994 18562 17006
rect 18510 16930 18562 16942
rect 19070 16994 19122 17006
rect 19070 16930 19122 16942
rect 24782 16994 24834 17006
rect 24782 16930 24834 16942
rect 27806 16994 27858 17006
rect 27806 16930 27858 16942
rect 2270 16882 2322 16894
rect 2270 16818 2322 16830
rect 3838 16882 3890 16894
rect 3838 16818 3890 16830
rect 4734 16882 4786 16894
rect 4734 16818 4786 16830
rect 7758 16882 7810 16894
rect 7758 16818 7810 16830
rect 8206 16882 8258 16894
rect 8206 16818 8258 16830
rect 10558 16882 10610 16894
rect 10558 16818 10610 16830
rect 11790 16882 11842 16894
rect 11790 16818 11842 16830
rect 14254 16882 14306 16894
rect 14254 16818 14306 16830
rect 14590 16882 14642 16894
rect 14590 16818 14642 16830
rect 14814 16882 14866 16894
rect 14814 16818 14866 16830
rect 14926 16882 14978 16894
rect 14926 16818 14978 16830
rect 15262 16882 15314 16894
rect 15822 16882 15874 16894
rect 15698 16879 15710 16882
rect 15262 16818 15314 16830
rect 15377 16833 15710 16879
rect 13694 16770 13746 16782
rect 15377 16770 15423 16833
rect 15698 16830 15710 16833
rect 15762 16830 15774 16882
rect 15822 16818 15874 16830
rect 16270 16882 16322 16894
rect 16270 16818 16322 16830
rect 16606 16882 16658 16894
rect 16606 16818 16658 16830
rect 19742 16882 19794 16894
rect 19742 16818 19794 16830
rect 20078 16882 20130 16894
rect 20078 16818 20130 16830
rect 21758 16882 21810 16894
rect 21758 16818 21810 16830
rect 26462 16882 26514 16894
rect 26462 16818 26514 16830
rect 20862 16770 20914 16782
rect 15362 16718 15374 16770
rect 15426 16718 15438 16770
rect 13694 16706 13746 16718
rect 20862 16706 20914 16718
rect 21422 16770 21474 16782
rect 21422 16706 21474 16718
rect 22206 16770 22258 16782
rect 22206 16706 22258 16718
rect 23102 16770 23154 16782
rect 23102 16706 23154 16718
rect 25678 16770 25730 16782
rect 25678 16706 25730 16718
rect 26126 16770 26178 16782
rect 26126 16706 26178 16718
rect 27022 16770 27074 16782
rect 27022 16706 27074 16718
rect 27470 16770 27522 16782
rect 27470 16706 27522 16718
rect 7646 16658 7698 16670
rect 7646 16594 7698 16606
rect 12686 16658 12738 16670
rect 12686 16594 12738 16606
rect 17838 16658 17890 16670
rect 20738 16606 20750 16658
rect 20802 16655 20814 16658
rect 21522 16655 21534 16658
rect 20802 16609 21534 16655
rect 20802 16606 20814 16609
rect 21522 16606 21534 16609
rect 21586 16606 21598 16658
rect 27010 16606 27022 16658
rect 27074 16655 27086 16658
rect 27682 16655 27694 16658
rect 27074 16609 27694 16655
rect 27074 16606 27086 16609
rect 27682 16606 27694 16609
rect 27746 16606 27758 16658
rect 17838 16594 17890 16606
rect 1344 16490 42560 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 42560 16490
rect 1344 16404 42560 16438
rect 2382 16322 2434 16334
rect 2382 16258 2434 16270
rect 5742 16322 5794 16334
rect 5742 16258 5794 16270
rect 6078 16322 6130 16334
rect 6078 16258 6130 16270
rect 12798 16322 12850 16334
rect 12798 16258 12850 16270
rect 18846 16322 18898 16334
rect 18846 16258 18898 16270
rect 20750 16322 20802 16334
rect 20750 16258 20802 16270
rect 4734 16210 4786 16222
rect 22766 16210 22818 16222
rect 10546 16158 10558 16210
rect 10610 16158 10622 16210
rect 13906 16158 13918 16210
rect 13970 16158 13982 16210
rect 4734 16146 4786 16158
rect 22766 16146 22818 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 29486 16210 29538 16222
rect 29486 16146 29538 16158
rect 29934 16210 29986 16222
rect 29934 16146 29986 16158
rect 1822 16098 1874 16110
rect 1822 16034 1874 16046
rect 2270 16098 2322 16110
rect 2270 16034 2322 16046
rect 3054 16098 3106 16110
rect 3054 16034 3106 16046
rect 3838 16098 3890 16110
rect 3838 16034 3890 16046
rect 6526 16098 6578 16110
rect 13694 16098 13746 16110
rect 7746 16046 7758 16098
rect 7810 16046 7822 16098
rect 6526 16034 6578 16046
rect 13694 16034 13746 16046
rect 17950 16098 18002 16110
rect 21534 16098 21586 16110
rect 20402 16046 20414 16098
rect 20466 16046 20478 16098
rect 21858 16046 21870 16098
rect 21922 16046 21934 16098
rect 17950 16034 18002 16046
rect 21534 16034 21586 16046
rect 4622 15986 4674 15998
rect 3950 15930 4002 15942
rect 2382 15874 2434 15886
rect 2382 15810 2434 15822
rect 3166 15874 3218 15886
rect 3166 15810 3218 15822
rect 3390 15874 3442 15886
rect 4622 15922 4674 15934
rect 4846 15986 4898 15998
rect 4846 15922 4898 15934
rect 5966 15986 6018 15998
rect 11118 15986 11170 15998
rect 8418 15934 8430 15986
rect 8482 15934 8494 15986
rect 5966 15922 6018 15934
rect 11118 15922 11170 15934
rect 11230 15986 11282 15998
rect 11230 15922 11282 15934
rect 11454 15986 11506 15998
rect 11454 15922 11506 15934
rect 11902 15986 11954 15998
rect 11902 15922 11954 15934
rect 12686 15986 12738 15998
rect 12686 15922 12738 15934
rect 12798 15986 12850 15998
rect 12798 15922 12850 15934
rect 14590 15986 14642 15998
rect 14590 15922 14642 15934
rect 14702 15986 14754 15998
rect 14702 15922 14754 15934
rect 15374 15986 15426 15998
rect 16494 15986 16546 15998
rect 15698 15934 15710 15986
rect 15762 15934 15774 15986
rect 15374 15922 15426 15934
rect 16494 15922 16546 15934
rect 17166 15986 17218 15998
rect 17166 15922 17218 15934
rect 17390 15986 17442 15998
rect 17390 15922 17442 15934
rect 18062 15986 18114 15998
rect 18062 15922 18114 15934
rect 18734 15986 18786 15998
rect 18734 15922 18786 15934
rect 19406 15986 19458 15998
rect 19406 15922 19458 15934
rect 20190 15986 20242 15998
rect 20190 15922 20242 15934
rect 20638 15986 20690 15998
rect 20638 15922 20690 15934
rect 3950 15866 4002 15878
rect 4174 15874 4226 15886
rect 3390 15810 3442 15822
rect 4174 15810 4226 15822
rect 6862 15874 6914 15886
rect 6862 15810 6914 15822
rect 7086 15874 7138 15886
rect 7086 15810 7138 15822
rect 7198 15874 7250 15886
rect 7198 15810 7250 15822
rect 12014 15874 12066 15886
rect 12014 15810 12066 15822
rect 12238 15874 12290 15886
rect 12238 15810 12290 15822
rect 13918 15874 13970 15886
rect 13918 15810 13970 15822
rect 14926 15874 14978 15886
rect 14926 15810 14978 15822
rect 16158 15874 16210 15886
rect 16158 15810 16210 15822
rect 16382 15874 16434 15886
rect 16382 15810 16434 15822
rect 17278 15874 17330 15886
rect 17278 15810 17330 15822
rect 18286 15874 18338 15886
rect 18286 15810 18338 15822
rect 19518 15874 19570 15886
rect 19518 15810 19570 15822
rect 19742 15874 19794 15886
rect 19742 15810 19794 15822
rect 22094 15874 22146 15886
rect 22094 15810 22146 15822
rect 22206 15874 22258 15886
rect 22206 15810 22258 15822
rect 22654 15874 22706 15886
rect 22654 15810 22706 15822
rect 23998 15874 24050 15886
rect 23998 15810 24050 15822
rect 24894 15874 24946 15886
rect 24894 15810 24946 15822
rect 25230 15874 25282 15886
rect 25230 15810 25282 15822
rect 26014 15874 26066 15886
rect 26014 15810 26066 15822
rect 26462 15874 26514 15886
rect 26462 15810 26514 15822
rect 26798 15874 26850 15886
rect 26798 15810 26850 15822
rect 27246 15874 27298 15886
rect 27246 15810 27298 15822
rect 27694 15874 27746 15886
rect 27694 15810 27746 15822
rect 28254 15874 28306 15886
rect 28254 15810 28306 15822
rect 28814 15874 28866 15886
rect 28814 15810 28866 15822
rect 1344 15706 42560 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 42560 15706
rect 1344 15620 42560 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 2270 15538 2322 15550
rect 2270 15474 2322 15486
rect 2830 15538 2882 15550
rect 2830 15474 2882 15486
rect 3054 15538 3106 15550
rect 3054 15474 3106 15486
rect 4398 15538 4450 15550
rect 4398 15474 4450 15486
rect 5182 15538 5234 15550
rect 5182 15474 5234 15486
rect 5406 15538 5458 15550
rect 5406 15474 5458 15486
rect 7310 15538 7362 15550
rect 7310 15474 7362 15486
rect 7534 15538 7586 15550
rect 7534 15474 7586 15486
rect 8318 15538 8370 15550
rect 8318 15474 8370 15486
rect 8430 15538 8482 15550
rect 8430 15474 8482 15486
rect 10334 15538 10386 15550
rect 10334 15474 10386 15486
rect 11902 15538 11954 15550
rect 11902 15474 11954 15486
rect 12574 15538 12626 15550
rect 12574 15474 12626 15486
rect 12798 15538 12850 15550
rect 12798 15474 12850 15486
rect 13582 15538 13634 15550
rect 13582 15474 13634 15486
rect 14142 15538 14194 15550
rect 14142 15474 14194 15486
rect 16942 15538 16994 15550
rect 16942 15474 16994 15486
rect 17838 15538 17890 15550
rect 17838 15474 17890 15486
rect 20750 15538 20802 15550
rect 20750 15474 20802 15486
rect 20862 15538 20914 15550
rect 20862 15474 20914 15486
rect 21310 15538 21362 15550
rect 21310 15474 21362 15486
rect 21534 15538 21586 15550
rect 21534 15474 21586 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 27134 15538 27186 15550
rect 27134 15474 27186 15486
rect 30718 15538 30770 15550
rect 30718 15474 30770 15486
rect 1934 15426 1986 15438
rect 1934 15362 1986 15374
rect 2718 15426 2770 15438
rect 2718 15362 2770 15374
rect 3502 15426 3554 15438
rect 3502 15362 3554 15374
rect 3614 15426 3666 15438
rect 3614 15362 3666 15374
rect 4286 15426 4338 15438
rect 4286 15362 4338 15374
rect 5070 15426 5122 15438
rect 5070 15362 5122 15374
rect 5854 15426 5906 15438
rect 5854 15362 5906 15374
rect 6302 15426 6354 15438
rect 6302 15362 6354 15374
rect 7086 15426 7138 15438
rect 7086 15362 7138 15374
rect 8094 15426 8146 15438
rect 8094 15362 8146 15374
rect 9998 15426 10050 15438
rect 9998 15362 10050 15374
rect 10110 15426 10162 15438
rect 10110 15362 10162 15374
rect 10894 15426 10946 15438
rect 10894 15362 10946 15374
rect 11678 15426 11730 15438
rect 11678 15362 11730 15374
rect 13358 15426 13410 15438
rect 13358 15362 13410 15374
rect 18622 15426 18674 15438
rect 18622 15362 18674 15374
rect 19742 15426 19794 15438
rect 19742 15362 19794 15374
rect 22766 15426 22818 15438
rect 22766 15362 22818 15374
rect 24446 15426 24498 15438
rect 24446 15362 24498 15374
rect 24558 15426 24610 15438
rect 24558 15362 24610 15374
rect 25678 15426 25730 15438
rect 25678 15362 25730 15374
rect 31166 15426 31218 15438
rect 31166 15362 31218 15374
rect 3838 15314 3890 15326
rect 3838 15250 3890 15262
rect 4622 15314 4674 15326
rect 4622 15250 4674 15262
rect 6078 15314 6130 15326
rect 6078 15250 6130 15262
rect 6414 15314 6466 15326
rect 6414 15250 6466 15262
rect 8542 15314 8594 15326
rect 10782 15314 10834 15326
rect 8754 15262 8766 15314
rect 8818 15262 8830 15314
rect 8542 15250 8594 15262
rect 10782 15250 10834 15262
rect 11118 15314 11170 15326
rect 11118 15250 11170 15262
rect 11566 15314 11618 15326
rect 11566 15250 11618 15262
rect 12238 15314 12290 15326
rect 12238 15250 12290 15262
rect 14590 15314 14642 15326
rect 14590 15250 14642 15262
rect 14926 15314 14978 15326
rect 14926 15250 14978 15262
rect 15262 15314 15314 15326
rect 15262 15250 15314 15262
rect 15710 15314 15762 15326
rect 15710 15250 15762 15262
rect 16158 15314 16210 15326
rect 16158 15250 16210 15262
rect 16270 15314 16322 15326
rect 16270 15250 16322 15262
rect 17614 15314 17666 15326
rect 17614 15250 17666 15262
rect 17950 15314 18002 15326
rect 17950 15250 18002 15262
rect 18510 15314 18562 15326
rect 18510 15250 18562 15262
rect 18734 15314 18786 15326
rect 18734 15250 18786 15262
rect 19182 15314 19234 15326
rect 19182 15250 19234 15262
rect 19630 15314 19682 15326
rect 21870 15314 21922 15326
rect 20290 15262 20302 15314
rect 20354 15262 20366 15314
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 19630 15250 19682 15262
rect 21870 15250 21922 15262
rect 22542 15314 22594 15326
rect 22542 15250 22594 15262
rect 23214 15314 23266 15326
rect 23214 15250 23266 15262
rect 28030 15314 28082 15326
rect 28030 15250 28082 15262
rect 29822 15314 29874 15326
rect 29822 15250 29874 15262
rect 12462 15202 12514 15214
rect 14814 15202 14866 15214
rect 7522 15150 7534 15202
rect 7586 15150 7598 15202
rect 13682 15150 13694 15202
rect 13746 15150 13758 15202
rect 12462 15138 12514 15150
rect 14814 15138 14866 15150
rect 15934 15202 15986 15214
rect 15934 15138 15986 15150
rect 22990 15202 23042 15214
rect 22990 15138 23042 15150
rect 23774 15202 23826 15214
rect 23774 15138 23826 15150
rect 25790 15202 25842 15214
rect 25790 15138 25842 15150
rect 26798 15202 26850 15214
rect 26798 15138 26850 15150
rect 27582 15202 27634 15214
rect 27582 15138 27634 15150
rect 28590 15202 28642 15214
rect 28590 15138 28642 15150
rect 29038 15202 29090 15214
rect 29038 15138 29090 15150
rect 29486 15202 29538 15214
rect 29486 15138 29538 15150
rect 30382 15202 30434 15214
rect 30382 15138 30434 15150
rect 31726 15202 31778 15214
rect 31726 15138 31778 15150
rect 32174 15202 32226 15214
rect 32174 15138 32226 15150
rect 32622 15202 32674 15214
rect 32622 15138 32674 15150
rect 21198 15090 21250 15102
rect 21198 15026 21250 15038
rect 23662 15090 23714 15102
rect 23662 15026 23714 15038
rect 24446 15090 24498 15102
rect 24446 15026 24498 15038
rect 1344 14922 42560 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 42560 14922
rect 1344 14836 42560 14870
rect 16270 14754 16322 14766
rect 16270 14690 16322 14702
rect 17390 14754 17442 14766
rect 17390 14690 17442 14702
rect 19406 14754 19458 14766
rect 31938 14702 31950 14754
rect 32002 14751 32014 14754
rect 33506 14751 33518 14754
rect 32002 14705 33518 14751
rect 32002 14702 32014 14705
rect 33506 14702 33518 14705
rect 33570 14702 33582 14754
rect 19406 14690 19458 14702
rect 12238 14642 12290 14654
rect 2146 14590 2158 14642
rect 2210 14590 2222 14642
rect 8754 14590 8766 14642
rect 8818 14590 8830 14642
rect 12238 14578 12290 14590
rect 14814 14642 14866 14654
rect 27470 14642 27522 14654
rect 23762 14590 23774 14642
rect 23826 14590 23838 14642
rect 25890 14590 25902 14642
rect 25954 14590 25966 14642
rect 14814 14578 14866 14590
rect 27470 14578 27522 14590
rect 28030 14642 28082 14654
rect 28030 14578 28082 14590
rect 3838 14530 3890 14542
rect 2370 14478 2382 14530
rect 2434 14478 2446 14530
rect 3838 14466 3890 14478
rect 6078 14530 6130 14542
rect 6078 14466 6130 14478
rect 8206 14530 8258 14542
rect 12686 14530 12738 14542
rect 11554 14478 11566 14530
rect 11618 14478 11630 14530
rect 8206 14466 8258 14478
rect 12686 14466 12738 14478
rect 13022 14530 13074 14542
rect 13022 14466 13074 14478
rect 14030 14530 14082 14542
rect 14030 14466 14082 14478
rect 15038 14530 15090 14542
rect 19518 14530 19570 14542
rect 27022 14530 27074 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 16818 14478 16830 14530
rect 16882 14478 16894 14530
rect 17042 14478 17054 14530
rect 17106 14478 17118 14530
rect 18386 14478 18398 14530
rect 18450 14478 18462 14530
rect 20066 14478 20078 14530
rect 20130 14478 20142 14530
rect 21634 14478 21646 14530
rect 21698 14478 21710 14530
rect 22978 14478 22990 14530
rect 23042 14478 23054 14530
rect 15038 14466 15090 14478
rect 19518 14466 19570 14478
rect 27022 14466 27074 14478
rect 3502 14418 3554 14430
rect 3502 14354 3554 14366
rect 4286 14418 4338 14430
rect 4286 14354 4338 14366
rect 7198 14418 7250 14430
rect 12798 14418 12850 14430
rect 10882 14366 10894 14418
rect 10946 14366 10958 14418
rect 7198 14354 7250 14366
rect 12798 14354 12850 14366
rect 14142 14418 14194 14430
rect 14142 14354 14194 14366
rect 15934 14418 15986 14430
rect 15934 14354 15986 14366
rect 18062 14418 18114 14430
rect 18062 14354 18114 14366
rect 20526 14418 20578 14430
rect 20526 14354 20578 14366
rect 21982 14418 22034 14430
rect 21982 14354 22034 14366
rect 33294 14418 33346 14430
rect 33294 14354 33346 14366
rect 2942 14306 2994 14318
rect 2942 14242 2994 14254
rect 3614 14306 3666 14318
rect 3614 14242 3666 14254
rect 4398 14306 4450 14318
rect 4398 14242 4450 14254
rect 5854 14306 5906 14318
rect 5854 14242 5906 14254
rect 5966 14306 6018 14318
rect 5966 14242 6018 14254
rect 6750 14306 6802 14318
rect 6750 14242 6802 14254
rect 7310 14306 7362 14318
rect 7310 14242 7362 14254
rect 7534 14306 7586 14318
rect 7534 14242 7586 14254
rect 7870 14306 7922 14318
rect 7870 14242 7922 14254
rect 8094 14306 8146 14318
rect 8094 14242 8146 14254
rect 14366 14306 14418 14318
rect 17278 14306 17330 14318
rect 15362 14254 15374 14306
rect 15426 14254 15438 14306
rect 14366 14242 14418 14254
rect 17278 14242 17330 14254
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 19406 14306 19458 14318
rect 19406 14242 19458 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 20638 14306 20690 14318
rect 20638 14242 20690 14254
rect 22094 14306 22146 14318
rect 22094 14242 22146 14254
rect 22206 14306 22258 14318
rect 22206 14242 22258 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 26462 14306 26514 14318
rect 26462 14242 26514 14254
rect 26686 14306 26738 14318
rect 26686 14242 26738 14254
rect 27582 14306 27634 14318
rect 27582 14242 27634 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 29598 14306 29650 14318
rect 29598 14242 29650 14254
rect 29934 14306 29986 14318
rect 29934 14242 29986 14254
rect 30382 14306 30434 14318
rect 30382 14242 30434 14254
rect 30942 14306 30994 14318
rect 30942 14242 30994 14254
rect 31614 14306 31666 14318
rect 31614 14242 31666 14254
rect 32062 14306 32114 14318
rect 32062 14242 32114 14254
rect 32398 14306 32450 14318
rect 32398 14242 32450 14254
rect 32846 14306 32898 14318
rect 32846 14242 32898 14254
rect 33854 14306 33906 14318
rect 33854 14242 33906 14254
rect 34302 14306 34354 14318
rect 34302 14242 34354 14254
rect 1344 14138 42560 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 42560 14138
rect 1344 14052 42560 14086
rect 8094 13970 8146 13982
rect 8094 13906 8146 13918
rect 8878 13970 8930 13982
rect 8878 13906 8930 13918
rect 10110 13970 10162 13982
rect 10110 13906 10162 13918
rect 10222 13970 10274 13982
rect 10222 13906 10274 13918
rect 10334 13970 10386 13982
rect 10334 13906 10386 13918
rect 11118 13970 11170 13982
rect 11118 13906 11170 13918
rect 11790 13970 11842 13982
rect 11790 13906 11842 13918
rect 12014 13970 12066 13982
rect 12014 13906 12066 13918
rect 12574 13970 12626 13982
rect 12574 13906 12626 13918
rect 13582 13970 13634 13982
rect 13582 13906 13634 13918
rect 14590 13970 14642 13982
rect 14590 13906 14642 13918
rect 17054 13970 17106 13982
rect 17054 13906 17106 13918
rect 19070 13970 19122 13982
rect 20190 13970 20242 13982
rect 19070 13906 19122 13918
rect 19630 13914 19682 13926
rect 6414 13858 6466 13870
rect 6414 13794 6466 13806
rect 7086 13858 7138 13870
rect 7086 13794 7138 13806
rect 7310 13858 7362 13870
rect 7310 13794 7362 13806
rect 8206 13858 8258 13870
rect 8206 13794 8258 13806
rect 8766 13858 8818 13870
rect 8766 13794 8818 13806
rect 12462 13858 12514 13870
rect 12462 13794 12514 13806
rect 12798 13858 12850 13870
rect 12798 13794 12850 13806
rect 13246 13858 13298 13870
rect 13246 13794 13298 13806
rect 13358 13858 13410 13870
rect 13358 13794 13410 13806
rect 14366 13858 14418 13870
rect 14366 13794 14418 13806
rect 14814 13858 14866 13870
rect 14814 13794 14866 13806
rect 15374 13858 15426 13870
rect 15374 13794 15426 13806
rect 15822 13858 15874 13870
rect 15822 13794 15874 13806
rect 16830 13858 16882 13870
rect 16830 13794 16882 13806
rect 18062 13858 18114 13870
rect 18062 13794 18114 13806
rect 18734 13858 18786 13870
rect 18734 13794 18786 13806
rect 18846 13858 18898 13870
rect 18846 13794 18898 13806
rect 19518 13858 19570 13870
rect 20190 13906 20242 13918
rect 20414 13970 20466 13982
rect 20414 13906 20466 13918
rect 21646 13970 21698 13982
rect 21646 13906 21698 13918
rect 21758 13970 21810 13982
rect 21758 13906 21810 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 28142 13970 28194 13982
rect 28142 13906 28194 13918
rect 32174 13970 32226 13982
rect 32174 13906 32226 13918
rect 19630 13850 19682 13862
rect 23326 13858 23378 13870
rect 19518 13794 19570 13806
rect 23326 13794 23378 13806
rect 24446 13858 24498 13870
rect 24446 13794 24498 13806
rect 27358 13858 27410 13870
rect 27358 13794 27410 13806
rect 6302 13746 6354 13758
rect 4834 13694 4846 13746
rect 4898 13694 4910 13746
rect 5506 13694 5518 13746
rect 5570 13694 5582 13746
rect 6302 13682 6354 13694
rect 7870 13746 7922 13758
rect 7870 13682 7922 13694
rect 9102 13746 9154 13758
rect 10446 13746 10498 13758
rect 9874 13694 9886 13746
rect 9938 13694 9950 13746
rect 9102 13682 9154 13694
rect 10446 13682 10498 13694
rect 11678 13746 11730 13758
rect 16718 13746 16770 13758
rect 15586 13694 15598 13746
rect 15650 13694 15662 13746
rect 11678 13682 11730 13694
rect 16718 13682 16770 13694
rect 17950 13746 18002 13758
rect 17950 13682 18002 13694
rect 19854 13746 19906 13758
rect 19854 13682 19906 13694
rect 20526 13746 20578 13758
rect 20526 13682 20578 13694
rect 21534 13746 21586 13758
rect 21534 13682 21586 13694
rect 22206 13746 22258 13758
rect 22206 13682 22258 13694
rect 23550 13746 23602 13758
rect 23550 13682 23602 13694
rect 26014 13746 26066 13758
rect 26014 13682 26066 13694
rect 26350 13746 26402 13758
rect 26350 13682 26402 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 27134 13746 27186 13758
rect 27134 13682 27186 13694
rect 27470 13746 27522 13758
rect 27470 13682 27522 13694
rect 27918 13746 27970 13758
rect 27918 13682 27970 13694
rect 28254 13746 28306 13758
rect 28254 13682 28306 13694
rect 29822 13746 29874 13758
rect 29822 13682 29874 13694
rect 20974 13634 21026 13646
rect 1922 13582 1934 13634
rect 1986 13582 1998 13634
rect 4050 13582 4062 13634
rect 4114 13582 4126 13634
rect 5730 13582 5742 13634
rect 5794 13582 5806 13634
rect 7410 13582 7422 13634
rect 7474 13582 7486 13634
rect 15474 13582 15486 13634
rect 15538 13582 15550 13634
rect 20974 13570 21026 13582
rect 22654 13634 22706 13646
rect 22654 13570 22706 13582
rect 22766 13634 22818 13646
rect 22766 13570 22818 13582
rect 25566 13634 25618 13646
rect 25566 13570 25618 13582
rect 26238 13634 26290 13646
rect 26238 13570 26290 13582
rect 28814 13634 28866 13646
rect 28814 13570 28866 13582
rect 29374 13634 29426 13646
rect 29374 13570 29426 13582
rect 30270 13634 30322 13646
rect 30270 13570 30322 13582
rect 30718 13634 30770 13646
rect 30718 13570 30770 13582
rect 31166 13634 31218 13646
rect 31166 13570 31218 13582
rect 31726 13634 31778 13646
rect 31726 13570 31778 13582
rect 32622 13634 32674 13646
rect 32622 13570 32674 13582
rect 33518 13634 33570 13646
rect 33518 13570 33570 13582
rect 34078 13634 34130 13646
rect 34078 13570 34130 13582
rect 34526 13634 34578 13646
rect 34526 13570 34578 13582
rect 34862 13634 34914 13646
rect 34862 13570 34914 13582
rect 35422 13634 35474 13646
rect 35422 13570 35474 13582
rect 35870 13634 35922 13646
rect 35870 13570 35922 13582
rect 6414 13522 6466 13534
rect 6414 13458 6466 13470
rect 14478 13522 14530 13534
rect 14478 13458 14530 13470
rect 18062 13522 18114 13534
rect 18062 13458 18114 13470
rect 23886 13522 23938 13534
rect 23886 13458 23938 13470
rect 24558 13522 24610 13534
rect 24558 13458 24610 13470
rect 28926 13522 28978 13534
rect 29586 13470 29598 13522
rect 29650 13519 29662 13522
rect 30258 13519 30270 13522
rect 29650 13473 30270 13519
rect 29650 13470 29662 13473
rect 30258 13470 30270 13473
rect 30322 13470 30334 13522
rect 33618 13470 33630 13522
rect 33682 13519 33694 13522
rect 34850 13519 34862 13522
rect 33682 13473 34862 13519
rect 33682 13470 33694 13473
rect 34850 13470 34862 13473
rect 34914 13470 34926 13522
rect 28926 13458 28978 13470
rect 1344 13354 42560 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 42560 13354
rect 1344 13268 42560 13302
rect 4622 13186 4674 13198
rect 4622 13122 4674 13134
rect 6078 13186 6130 13198
rect 6078 13122 6130 13134
rect 14366 13186 14418 13198
rect 14366 13122 14418 13134
rect 14926 13186 14978 13198
rect 14926 13122 14978 13134
rect 25566 13186 25618 13198
rect 25566 13122 25618 13134
rect 27470 13186 27522 13198
rect 33506 13134 33518 13186
rect 33570 13183 33582 13186
rect 35970 13183 35982 13186
rect 33570 13137 35982 13183
rect 33570 13134 33582 13137
rect 35970 13134 35982 13137
rect 36034 13134 36046 13186
rect 27470 13122 27522 13134
rect 3950 13074 4002 13086
rect 3950 13010 4002 13022
rect 7310 13074 7362 13086
rect 7310 13010 7362 13022
rect 8206 13074 8258 13086
rect 24446 13074 24498 13086
rect 9650 13022 9662 13074
rect 9714 13022 9726 13074
rect 8206 13010 8258 13022
rect 24446 13010 24498 13022
rect 33742 13074 33794 13086
rect 33742 13010 33794 13022
rect 3166 12962 3218 12974
rect 5966 12962 6018 12974
rect 2034 12910 2046 12962
rect 2098 12910 2110 12962
rect 5730 12910 5742 12962
rect 5794 12910 5806 12962
rect 3166 12898 3218 12910
rect 5966 12898 6018 12910
rect 8430 12962 8482 12974
rect 14590 12962 14642 12974
rect 12562 12910 12574 12962
rect 12626 12910 12638 12962
rect 8430 12898 8482 12910
rect 14590 12898 14642 12910
rect 14814 12962 14866 12974
rect 14814 12898 14866 12910
rect 15710 12962 15762 12974
rect 15710 12898 15762 12910
rect 15822 12962 15874 12974
rect 15822 12898 15874 12910
rect 16270 12962 16322 12974
rect 16270 12898 16322 12910
rect 16606 12962 16658 12974
rect 16606 12898 16658 12910
rect 18958 12962 19010 12974
rect 18958 12898 19010 12910
rect 19294 12962 19346 12974
rect 19294 12898 19346 12910
rect 20078 12962 20130 12974
rect 20078 12898 20130 12910
rect 20414 12962 20466 12974
rect 24670 12962 24722 12974
rect 23314 12910 23326 12962
rect 23378 12910 23390 12962
rect 23538 12910 23550 12962
rect 23602 12910 23614 12962
rect 20414 12898 20466 12910
rect 24670 12898 24722 12910
rect 26238 12962 26290 12974
rect 26238 12898 26290 12910
rect 26462 12962 26514 12974
rect 26462 12898 26514 12910
rect 26910 12962 26962 12974
rect 26910 12898 26962 12910
rect 32846 12962 32898 12974
rect 32846 12898 32898 12910
rect 4062 12850 4114 12862
rect 2258 12798 2270 12850
rect 2322 12798 2334 12850
rect 4062 12786 4114 12798
rect 6974 12850 7026 12862
rect 13694 12850 13746 12862
rect 11778 12798 11790 12850
rect 11842 12798 11854 12850
rect 6974 12786 7026 12798
rect 13694 12786 13746 12798
rect 14254 12850 14306 12862
rect 14254 12786 14306 12798
rect 17166 12850 17218 12862
rect 17726 12850 17778 12862
rect 17378 12798 17390 12850
rect 17442 12847 17454 12850
rect 17602 12847 17614 12850
rect 17442 12801 17614 12847
rect 17442 12798 17454 12801
rect 17602 12798 17614 12801
rect 17666 12798 17678 12850
rect 17166 12786 17218 12798
rect 17726 12786 17778 12798
rect 19742 12850 19794 12862
rect 19742 12786 19794 12798
rect 21870 12850 21922 12862
rect 21870 12786 21922 12798
rect 22542 12850 22594 12862
rect 22542 12786 22594 12798
rect 22654 12850 22706 12862
rect 22654 12786 22706 12798
rect 23774 12850 23826 12862
rect 23774 12786 23826 12798
rect 25678 12850 25730 12862
rect 25678 12786 25730 12798
rect 27358 12850 27410 12862
rect 27358 12786 27410 12798
rect 27470 12850 27522 12862
rect 27470 12786 27522 12798
rect 28254 12850 28306 12862
rect 28254 12786 28306 12798
rect 28366 12850 28418 12862
rect 28366 12786 28418 12798
rect 29598 12850 29650 12862
rect 29598 12786 29650 12798
rect 30270 12850 30322 12862
rect 30270 12786 30322 12798
rect 30942 12850 30994 12862
rect 30942 12786 30994 12798
rect 31726 12850 31778 12862
rect 31726 12786 31778 12798
rect 32286 12850 32338 12862
rect 32286 12786 32338 12798
rect 35534 12850 35586 12862
rect 35534 12786 35586 12798
rect 3054 12738 3106 12750
rect 3054 12674 3106 12686
rect 3838 12738 3890 12750
rect 3838 12674 3890 12686
rect 4734 12738 4786 12750
rect 4734 12674 4786 12686
rect 4846 12738 4898 12750
rect 4846 12674 4898 12686
rect 7198 12738 7250 12750
rect 7198 12674 7250 12686
rect 7422 12738 7474 12750
rect 7422 12674 7474 12686
rect 7534 12738 7586 12750
rect 15934 12738 15986 12750
rect 8754 12686 8766 12738
rect 8818 12686 8830 12738
rect 7534 12674 7586 12686
rect 15934 12674 15986 12686
rect 16942 12738 16994 12750
rect 16942 12674 16994 12686
rect 17278 12738 17330 12750
rect 17278 12674 17330 12686
rect 17838 12738 17890 12750
rect 17838 12674 17890 12686
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 20190 12738 20242 12750
rect 20190 12674 20242 12686
rect 20862 12738 20914 12750
rect 20862 12674 20914 12686
rect 21534 12738 21586 12750
rect 21534 12674 21586 12686
rect 21758 12738 21810 12750
rect 21758 12674 21810 12686
rect 22318 12738 22370 12750
rect 22318 12674 22370 12686
rect 23886 12738 23938 12750
rect 26350 12738 26402 12750
rect 24994 12686 25006 12738
rect 25058 12686 25070 12738
rect 23886 12674 23938 12686
rect 26350 12674 26402 12686
rect 28030 12738 28082 12750
rect 28030 12674 28082 12686
rect 28814 12738 28866 12750
rect 28814 12674 28866 12686
rect 29710 12738 29762 12750
rect 29710 12674 29762 12686
rect 30382 12738 30434 12750
rect 30382 12674 30434 12686
rect 31054 12738 31106 12750
rect 31054 12674 31106 12686
rect 31614 12738 31666 12750
rect 31614 12674 31666 12686
rect 32398 12738 32450 12750
rect 32398 12674 32450 12686
rect 33294 12738 33346 12750
rect 33294 12674 33346 12686
rect 34190 12738 34242 12750
rect 34190 12674 34242 12686
rect 34750 12738 34802 12750
rect 34750 12674 34802 12686
rect 35086 12738 35138 12750
rect 35086 12674 35138 12686
rect 35982 12738 36034 12750
rect 35982 12674 36034 12686
rect 36430 12738 36482 12750
rect 36430 12674 36482 12686
rect 37438 12738 37490 12750
rect 37438 12674 37490 12686
rect 37886 12738 37938 12750
rect 37886 12674 37938 12686
rect 1344 12570 42560 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 42560 12570
rect 1344 12484 42560 12518
rect 1934 12402 1986 12414
rect 1934 12338 1986 12350
rect 2606 12402 2658 12414
rect 2606 12338 2658 12350
rect 3726 12402 3778 12414
rect 3726 12338 3778 12350
rect 4622 12402 4674 12414
rect 4622 12338 4674 12350
rect 5406 12402 5458 12414
rect 5406 12338 5458 12350
rect 6750 12402 6802 12414
rect 6750 12338 6802 12350
rect 6974 12402 7026 12414
rect 6974 12338 7026 12350
rect 8206 12402 8258 12414
rect 8206 12338 8258 12350
rect 8430 12402 8482 12414
rect 8430 12338 8482 12350
rect 9102 12402 9154 12414
rect 9102 12338 9154 12350
rect 17614 12402 17666 12414
rect 17614 12338 17666 12350
rect 18846 12402 18898 12414
rect 18846 12338 18898 12350
rect 23214 12402 23266 12414
rect 25566 12402 25618 12414
rect 24210 12350 24222 12402
rect 24274 12350 24286 12402
rect 23214 12338 23266 12350
rect 25566 12338 25618 12350
rect 25790 12402 25842 12414
rect 25790 12338 25842 12350
rect 33518 12402 33570 12414
rect 33518 12338 33570 12350
rect 34862 12402 34914 12414
rect 34862 12338 34914 12350
rect 36542 12402 36594 12414
rect 36542 12338 36594 12350
rect 40462 12402 40514 12414
rect 40462 12338 40514 12350
rect 41470 12402 41522 12414
rect 41470 12338 41522 12350
rect 42030 12402 42082 12414
rect 42030 12338 42082 12350
rect 1822 12290 1874 12302
rect 1822 12226 1874 12238
rect 2494 12290 2546 12302
rect 2494 12226 2546 12238
rect 3950 12290 4002 12302
rect 3950 12226 4002 12238
rect 4510 12290 4562 12302
rect 4510 12226 4562 12238
rect 5182 12290 5234 12302
rect 5182 12226 5234 12238
rect 5630 12290 5682 12302
rect 5630 12226 5682 12238
rect 11006 12290 11058 12302
rect 11006 12226 11058 12238
rect 17838 12290 17890 12302
rect 17838 12226 17890 12238
rect 17950 12290 18002 12302
rect 17950 12226 18002 12238
rect 18622 12290 18674 12302
rect 23102 12290 23154 12302
rect 20290 12238 20302 12290
rect 20354 12238 20366 12290
rect 18622 12226 18674 12238
rect 23102 12226 23154 12238
rect 23662 12290 23714 12302
rect 23662 12226 23714 12238
rect 25902 12290 25954 12302
rect 30270 12290 30322 12302
rect 27458 12238 27470 12290
rect 27522 12238 27534 12290
rect 25902 12226 25954 12238
rect 30270 12226 30322 12238
rect 32734 12290 32786 12302
rect 32734 12226 32786 12238
rect 33966 12290 34018 12302
rect 33966 12226 34018 12238
rect 3502 12178 3554 12190
rect 2818 12126 2830 12178
rect 2882 12126 2894 12178
rect 3502 12114 3554 12126
rect 3726 12178 3778 12190
rect 3726 12114 3778 12126
rect 7422 12178 7474 12190
rect 9774 12178 9826 12190
rect 18510 12178 18562 12190
rect 23326 12178 23378 12190
rect 7970 12126 7982 12178
rect 8034 12126 8046 12178
rect 16706 12126 16718 12178
rect 16770 12126 16782 12178
rect 19618 12126 19630 12178
rect 19682 12126 19694 12178
rect 7422 12114 7474 12126
rect 9774 12114 9826 12126
rect 18510 12114 18562 12126
rect 23326 12114 23378 12126
rect 23438 12178 23490 12190
rect 23438 12114 23490 12126
rect 24558 12178 24610 12190
rect 30158 12178 30210 12190
rect 26674 12126 26686 12178
rect 26738 12126 26750 12178
rect 24558 12114 24610 12126
rect 30158 12114 30210 12126
rect 32846 12178 32898 12190
rect 32846 12114 32898 12126
rect 6302 12066 6354 12078
rect 6302 12002 6354 12014
rect 6862 12066 6914 12078
rect 6862 12002 6914 12014
rect 8094 12066 8146 12078
rect 24782 12066 24834 12078
rect 30942 12066 30994 12078
rect 10210 12014 10222 12066
rect 10274 12014 10286 12066
rect 14578 12014 14590 12066
rect 14642 12014 14654 12066
rect 22418 12014 22430 12066
rect 22482 12014 22494 12066
rect 29586 12014 29598 12066
rect 29650 12014 29662 12066
rect 8094 12002 8146 12014
rect 24782 12002 24834 12014
rect 30942 12002 30994 12014
rect 31614 12066 31666 12078
rect 31614 12002 31666 12014
rect 32062 12066 32114 12078
rect 32062 12002 32114 12014
rect 34414 12066 34466 12078
rect 34414 12002 34466 12014
rect 35646 12066 35698 12078
rect 35646 12002 35698 12014
rect 36094 12066 36146 12078
rect 36094 12002 36146 12014
rect 36990 12066 37042 12078
rect 36990 12002 37042 12014
rect 37886 12066 37938 12078
rect 37886 12002 37938 12014
rect 37998 12066 38050 12078
rect 37998 12002 38050 12014
rect 38558 12066 38610 12078
rect 38558 12002 38610 12014
rect 38894 12066 38946 12078
rect 38894 12002 38946 12014
rect 39566 12066 39618 12078
rect 39566 12002 39618 12014
rect 5742 11954 5794 11966
rect 5742 11890 5794 11902
rect 10894 11954 10946 11966
rect 10894 11890 10946 11902
rect 30830 11954 30882 11966
rect 30830 11890 30882 11902
rect 31502 11954 31554 11966
rect 31502 11890 31554 11902
rect 32734 11954 32786 11966
rect 35534 11954 35586 11966
rect 33506 11902 33518 11954
rect 33570 11951 33582 11954
rect 33842 11951 33854 11954
rect 33570 11905 33854 11951
rect 33570 11902 33582 11905
rect 33842 11902 33854 11905
rect 33906 11951 33918 11954
rect 34402 11951 34414 11954
rect 33906 11905 34414 11951
rect 33906 11902 33918 11905
rect 34402 11902 34414 11905
rect 34466 11902 34478 11954
rect 32734 11890 32786 11902
rect 35534 11890 35586 11902
rect 1344 11786 42560 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 42560 11786
rect 1344 11700 42560 11734
rect 9326 11618 9378 11630
rect 9326 11554 9378 11566
rect 10782 11618 10834 11630
rect 10782 11554 10834 11566
rect 15934 11618 15986 11630
rect 40786 11566 40798 11618
rect 40850 11615 40862 11618
rect 41682 11615 41694 11618
rect 40850 11569 41694 11615
rect 40850 11566 40862 11569
rect 41682 11566 41694 11569
rect 41746 11566 41758 11618
rect 15934 11554 15986 11566
rect 7310 11506 7362 11518
rect 1810 11454 1822 11506
rect 1874 11454 1886 11506
rect 7310 11442 7362 11454
rect 8990 11506 9042 11518
rect 8990 11442 9042 11454
rect 12574 11506 12626 11518
rect 18174 11506 18226 11518
rect 27918 11506 27970 11518
rect 41694 11506 41746 11518
rect 14018 11454 14030 11506
rect 14082 11454 14094 11506
rect 21858 11454 21870 11506
rect 21922 11454 21934 11506
rect 36754 11454 36766 11506
rect 36818 11454 36830 11506
rect 12574 11442 12626 11454
rect 18174 11442 18226 11454
rect 27918 11442 27970 11454
rect 41694 11442 41746 11454
rect 6078 11394 6130 11406
rect 4722 11342 4734 11394
rect 4786 11342 4798 11394
rect 5730 11342 5742 11394
rect 5794 11342 5806 11394
rect 6078 11330 6130 11342
rect 6190 11394 6242 11406
rect 6190 11330 6242 11342
rect 6414 11394 6466 11406
rect 6414 11330 6466 11342
rect 6638 11394 6690 11406
rect 6638 11330 6690 11342
rect 7086 11394 7138 11406
rect 7086 11330 7138 11342
rect 7534 11394 7586 11406
rect 7534 11330 7586 11342
rect 8878 11394 8930 11406
rect 8878 11330 8930 11342
rect 9102 11394 9154 11406
rect 10222 11394 10274 11406
rect 11006 11394 11058 11406
rect 9538 11342 9550 11394
rect 9602 11342 9614 11394
rect 9762 11342 9774 11394
rect 9826 11342 9838 11394
rect 10546 11342 10558 11394
rect 10610 11342 10622 11394
rect 9102 11330 9154 11342
rect 10222 11330 10274 11342
rect 11006 11330 11058 11342
rect 11230 11394 11282 11406
rect 12686 11394 12738 11406
rect 17390 11394 17442 11406
rect 22206 11394 22258 11406
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 12898 11342 12910 11394
rect 12962 11342 12974 11394
rect 19394 11342 19406 11394
rect 19458 11342 19470 11394
rect 20402 11342 20414 11394
rect 20466 11342 20478 11394
rect 21634 11342 21646 11394
rect 21698 11342 21710 11394
rect 11230 11330 11282 11342
rect 12686 11330 12738 11342
rect 17390 11330 17442 11342
rect 22206 11330 22258 11342
rect 23550 11394 23602 11406
rect 23550 11330 23602 11342
rect 23886 11394 23938 11406
rect 23886 11330 23938 11342
rect 23998 11394 24050 11406
rect 23998 11330 24050 11342
rect 24558 11394 24610 11406
rect 24558 11330 24610 11342
rect 25678 11394 25730 11406
rect 25678 11330 25730 11342
rect 26014 11394 26066 11406
rect 26014 11330 26066 11342
rect 26686 11394 26738 11406
rect 26686 11330 26738 11342
rect 28366 11394 28418 11406
rect 28366 11330 28418 11342
rect 28702 11394 28754 11406
rect 28702 11330 28754 11342
rect 29934 11394 29986 11406
rect 29934 11330 29986 11342
rect 30606 11394 30658 11406
rect 30606 11330 30658 11342
rect 31726 11394 31778 11406
rect 31726 11330 31778 11342
rect 33182 11394 33234 11406
rect 37662 11394 37714 11406
rect 33842 11342 33854 11394
rect 33906 11342 33918 11394
rect 33182 11330 33234 11342
rect 37662 11330 37714 11342
rect 37886 11394 37938 11406
rect 37886 11330 37938 11342
rect 37998 11394 38050 11406
rect 39006 11394 39058 11406
rect 38658 11342 38670 11394
rect 38722 11342 38734 11394
rect 37998 11330 38050 11342
rect 39006 11330 39058 11342
rect 39230 11394 39282 11406
rect 39230 11330 39282 11342
rect 7758 11282 7810 11294
rect 3938 11230 3950 11282
rect 4002 11230 4014 11282
rect 7758 11218 7810 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 14702 11282 14754 11294
rect 14702 11218 14754 11230
rect 16158 11282 16210 11294
rect 16158 11218 16210 11230
rect 17502 11282 17554 11294
rect 17502 11218 17554 11230
rect 18622 11282 18674 11294
rect 18622 11218 18674 11230
rect 24894 11282 24946 11294
rect 24894 11218 24946 11230
rect 25790 11282 25842 11294
rect 25790 11218 25842 11230
rect 27470 11282 27522 11294
rect 27470 11218 27522 11230
rect 29598 11282 29650 11294
rect 29598 11218 29650 11230
rect 31054 11282 31106 11294
rect 31054 11218 31106 11230
rect 31838 11282 31890 11294
rect 31838 11218 31890 11230
rect 32510 11282 32562 11294
rect 32510 11218 32562 11230
rect 32622 11282 32674 11294
rect 37550 11282 37602 11294
rect 34626 11230 34638 11282
rect 34690 11230 34702 11282
rect 32622 11218 32674 11230
rect 37550 11218 37602 11230
rect 8318 11170 8370 11182
rect 11678 11170 11730 11182
rect 6066 11118 6078 11170
rect 6130 11118 6142 11170
rect 10658 11118 10670 11170
rect 10722 11118 10734 11170
rect 8318 11106 8370 11118
rect 11678 11106 11730 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 14814 11170 14866 11182
rect 17166 11170 17218 11182
rect 15586 11118 15598 11170
rect 15650 11118 15662 11170
rect 14814 11106 14866 11118
rect 17166 11106 17218 11118
rect 17614 11170 17666 11182
rect 17614 11106 17666 11118
rect 18734 11170 18786 11182
rect 18734 11106 18786 11118
rect 18958 11170 19010 11182
rect 18958 11106 19010 11118
rect 19630 11170 19682 11182
rect 19630 11106 19682 11118
rect 19854 11170 19906 11182
rect 19854 11106 19906 11118
rect 19966 11170 20018 11182
rect 19966 11106 20018 11118
rect 20638 11170 20690 11182
rect 20638 11106 20690 11118
rect 20862 11170 20914 11182
rect 20862 11106 20914 11118
rect 20974 11170 21026 11182
rect 20974 11106 21026 11118
rect 21870 11170 21922 11182
rect 21870 11106 21922 11118
rect 22094 11170 22146 11182
rect 22094 11106 22146 11118
rect 22766 11170 22818 11182
rect 22766 11106 22818 11118
rect 23662 11170 23714 11182
rect 23662 11106 23714 11118
rect 23774 11170 23826 11182
rect 23774 11106 23826 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 26350 11170 26402 11182
rect 26350 11106 26402 11118
rect 26574 11170 26626 11182
rect 26574 11106 26626 11118
rect 27134 11170 27186 11182
rect 27134 11106 27186 11118
rect 27358 11170 27410 11182
rect 27358 11106 27410 11118
rect 28590 11170 28642 11182
rect 28590 11106 28642 11118
rect 29710 11170 29762 11182
rect 29710 11106 29762 11118
rect 30270 11170 30322 11182
rect 30270 11106 30322 11118
rect 30494 11170 30546 11182
rect 30494 11106 30546 11118
rect 32062 11170 32114 11182
rect 32062 11106 32114 11118
rect 32846 11170 32898 11182
rect 32846 11106 32898 11118
rect 39678 11170 39730 11182
rect 39678 11106 39730 11118
rect 40350 11170 40402 11182
rect 40350 11106 40402 11118
rect 40798 11170 40850 11182
rect 40798 11106 40850 11118
rect 41246 11170 41298 11182
rect 41246 11106 41298 11118
rect 1344 11002 42560 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 42560 11002
rect 1344 10916 42560 10950
rect 4174 10834 4226 10846
rect 4174 10770 4226 10782
rect 4286 10834 4338 10846
rect 4286 10770 4338 10782
rect 4398 10834 4450 10846
rect 4398 10770 4450 10782
rect 4510 10834 4562 10846
rect 4510 10770 4562 10782
rect 6638 10834 6690 10846
rect 6638 10770 6690 10782
rect 7422 10834 7474 10846
rect 7422 10770 7474 10782
rect 8430 10834 8482 10846
rect 8430 10770 8482 10782
rect 9662 10834 9714 10846
rect 9662 10770 9714 10782
rect 15486 10834 15538 10846
rect 15486 10770 15538 10782
rect 15710 10834 15762 10846
rect 15710 10770 15762 10782
rect 16270 10834 16322 10846
rect 16270 10770 16322 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 32846 10834 32898 10846
rect 32846 10770 32898 10782
rect 34862 10834 34914 10846
rect 34862 10770 34914 10782
rect 35422 10834 35474 10846
rect 35422 10770 35474 10782
rect 36094 10834 36146 10846
rect 36094 10770 36146 10782
rect 38222 10834 38274 10846
rect 38222 10770 38274 10782
rect 40574 10834 40626 10846
rect 40574 10770 40626 10782
rect 41470 10834 41522 10846
rect 41470 10770 41522 10782
rect 5182 10722 5234 10734
rect 1922 10670 1934 10722
rect 1986 10670 1998 10722
rect 5182 10658 5234 10670
rect 5630 10722 5682 10734
rect 5630 10658 5682 10670
rect 7198 10722 7250 10734
rect 7198 10658 7250 10670
rect 7534 10722 7586 10734
rect 7534 10658 7586 10670
rect 10670 10722 10722 10734
rect 10670 10658 10722 10670
rect 15374 10722 15426 10734
rect 15374 10658 15426 10670
rect 16494 10722 16546 10734
rect 16494 10658 16546 10670
rect 17054 10722 17106 10734
rect 17054 10658 17106 10670
rect 17838 10722 17890 10734
rect 17838 10658 17890 10670
rect 33966 10722 34018 10734
rect 33966 10658 34018 10670
rect 36206 10722 36258 10734
rect 36206 10658 36258 10670
rect 36878 10722 36930 10734
rect 36878 10658 36930 10670
rect 7758 10610 7810 10622
rect 3938 10558 3950 10610
rect 4002 10558 4014 10610
rect 5394 10558 5406 10610
rect 5458 10558 5470 10610
rect 6178 10558 6190 10610
rect 6242 10558 6254 10610
rect 6402 10558 6414 10610
rect 6466 10558 6478 10610
rect 7758 10546 7810 10558
rect 9774 10610 9826 10622
rect 9774 10546 9826 10558
rect 9998 10610 10050 10622
rect 9998 10546 10050 10558
rect 10334 10610 10386 10622
rect 10334 10546 10386 10558
rect 11230 10610 11282 10622
rect 17950 10610 18002 10622
rect 24222 10610 24274 10622
rect 14690 10558 14702 10610
rect 14754 10558 14766 10610
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 11230 10546 11282 10558
rect 17950 10546 18002 10558
rect 24222 10546 24274 10558
rect 24558 10610 24610 10622
rect 24558 10546 24610 10558
rect 24894 10610 24946 10622
rect 33518 10610 33570 10622
rect 26002 10558 26014 10610
rect 26066 10558 26078 10610
rect 29586 10558 29598 10610
rect 29650 10558 29662 10610
rect 24894 10546 24946 10558
rect 33518 10546 33570 10558
rect 34190 10610 34242 10622
rect 34190 10546 34242 10558
rect 34750 10610 34802 10622
rect 34750 10546 34802 10558
rect 35870 10610 35922 10622
rect 35870 10546 35922 10558
rect 36990 10610 37042 10622
rect 36990 10546 37042 10558
rect 37998 10610 38050 10622
rect 37998 10546 38050 10558
rect 40126 10610 40178 10622
rect 40126 10546 40178 10558
rect 6750 10498 6802 10510
rect 3266 10446 3278 10498
rect 3330 10446 3342 10498
rect 6750 10434 6802 10446
rect 8990 10498 9042 10510
rect 24446 10498 24498 10510
rect 33742 10498 33794 10510
rect 11890 10446 11902 10498
rect 11954 10446 11966 10498
rect 14018 10446 14030 10498
rect 14082 10446 14094 10498
rect 20514 10446 20526 10498
rect 20578 10446 20590 10498
rect 26786 10446 26798 10498
rect 26850 10446 26862 10498
rect 28914 10446 28926 10498
rect 28978 10446 28990 10498
rect 30258 10446 30270 10498
rect 30322 10446 30334 10498
rect 32386 10446 32398 10498
rect 32450 10446 32462 10498
rect 8990 10434 9042 10446
rect 24446 10434 24498 10446
rect 33742 10434 33794 10446
rect 37438 10498 37490 10510
rect 38782 10498 38834 10510
rect 38210 10446 38222 10498
rect 38274 10446 38286 10498
rect 37438 10434 37490 10446
rect 38782 10434 38834 10446
rect 39230 10498 39282 10510
rect 39230 10434 39282 10446
rect 39678 10498 39730 10510
rect 39678 10434 39730 10446
rect 41918 10498 41970 10510
rect 41918 10434 41970 10446
rect 5294 10386 5346 10398
rect 5294 10322 5346 10334
rect 10222 10386 10274 10398
rect 10222 10322 10274 10334
rect 11342 10386 11394 10398
rect 11342 10322 11394 10334
rect 34862 10386 34914 10398
rect 34862 10322 34914 10334
rect 36878 10386 36930 10398
rect 36878 10322 36930 10334
rect 1344 10218 42560 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 42560 10218
rect 1344 10132 42560 10166
rect 4958 10050 5010 10062
rect 4958 9986 5010 9998
rect 7310 10050 7362 10062
rect 7310 9986 7362 9998
rect 10110 10050 10162 10062
rect 10110 9986 10162 9998
rect 17166 10050 17218 10062
rect 17166 9986 17218 9998
rect 27358 10050 27410 10062
rect 27358 9986 27410 9998
rect 27806 10050 27858 10062
rect 27806 9986 27858 9998
rect 2718 9938 2770 9950
rect 4846 9938 4898 9950
rect 2146 9886 2158 9938
rect 2210 9886 2222 9938
rect 3042 9886 3054 9938
rect 3106 9886 3118 9938
rect 2718 9874 2770 9886
rect 4846 9874 4898 9886
rect 6414 9938 6466 9950
rect 6414 9874 6466 9886
rect 14030 9938 14082 9950
rect 18510 9938 18562 9950
rect 16034 9886 16046 9938
rect 16098 9886 16110 9938
rect 14030 9874 14082 9886
rect 18510 9874 18562 9886
rect 21870 9938 21922 9950
rect 21870 9874 21922 9886
rect 22878 9938 22930 9950
rect 26686 9938 26738 9950
rect 24098 9886 24110 9938
rect 24162 9886 24174 9938
rect 26226 9886 26238 9938
rect 26290 9886 26302 9938
rect 22878 9874 22930 9886
rect 26686 9874 26738 9886
rect 27470 9938 27522 9950
rect 27470 9874 27522 9886
rect 27694 9938 27746 9950
rect 30158 9938 30210 9950
rect 37662 9938 37714 9950
rect 40574 9938 40626 9950
rect 28466 9886 28478 9938
rect 28530 9886 28542 9938
rect 33282 9886 33294 9938
rect 33346 9886 33358 9938
rect 35410 9886 35422 9938
rect 35474 9886 35486 9938
rect 38658 9886 38670 9938
rect 38722 9886 38734 9938
rect 27694 9874 27746 9886
rect 30158 9874 30210 9886
rect 37662 9874 37714 9886
rect 40574 9874 40626 9886
rect 41470 9938 41522 9950
rect 41470 9874 41522 9886
rect 41918 9938 41970 9950
rect 41918 9874 41970 9886
rect 3838 9826 3890 9838
rect 3838 9762 3890 9774
rect 4062 9826 4114 9838
rect 4062 9762 4114 9774
rect 6190 9826 6242 9838
rect 6190 9762 6242 9774
rect 7646 9826 7698 9838
rect 7646 9762 7698 9774
rect 9774 9826 9826 9838
rect 9774 9762 9826 9774
rect 10222 9826 10274 9838
rect 10222 9762 10274 9774
rect 11566 9826 11618 9838
rect 13918 9826 13970 9838
rect 13682 9774 13694 9826
rect 13746 9774 13758 9826
rect 11566 9762 11618 9774
rect 13918 9762 13970 9774
rect 14142 9826 14194 9838
rect 17726 9826 17778 9838
rect 14354 9774 14366 9826
rect 14418 9774 14430 9826
rect 16146 9774 16158 9826
rect 16210 9774 16222 9826
rect 14142 9762 14194 9774
rect 17726 9762 17778 9774
rect 18622 9826 18674 9838
rect 18622 9762 18674 9774
rect 18846 9826 18898 9838
rect 18846 9762 18898 9774
rect 20638 9826 20690 9838
rect 20638 9762 20690 9774
rect 20862 9826 20914 9838
rect 20862 9762 20914 9774
rect 22430 9826 22482 9838
rect 29822 9826 29874 9838
rect 23426 9774 23438 9826
rect 23490 9774 23502 9826
rect 22430 9762 22482 9774
rect 29822 9762 29874 9774
rect 30046 9826 30098 9838
rect 30046 9762 30098 9774
rect 30382 9826 30434 9838
rect 30382 9762 30434 9774
rect 31838 9826 31890 9838
rect 36206 9826 36258 9838
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 31838 9762 31890 9774
rect 36206 9762 36258 9774
rect 37886 9826 37938 9838
rect 40126 9826 40178 9838
rect 38098 9774 38110 9826
rect 38162 9774 38174 9826
rect 37886 9762 37938 9774
rect 40126 9762 40178 9774
rect 41022 9826 41074 9838
rect 41022 9762 41074 9774
rect 1822 9714 1874 9726
rect 1822 9650 1874 9662
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 3614 9714 3666 9726
rect 3614 9650 3666 9662
rect 5742 9714 5794 9726
rect 6638 9714 6690 9726
rect 5954 9662 5966 9714
rect 6018 9662 6030 9714
rect 5742 9650 5794 9662
rect 6638 9650 6690 9662
rect 7870 9714 7922 9726
rect 7870 9650 7922 9662
rect 8990 9714 9042 9726
rect 8990 9650 9042 9662
rect 9550 9714 9602 9726
rect 9550 9650 9602 9662
rect 10782 9714 10834 9726
rect 10782 9650 10834 9662
rect 12126 9714 12178 9726
rect 12126 9650 12178 9662
rect 12686 9714 12738 9726
rect 12686 9650 12738 9662
rect 12798 9714 12850 9726
rect 12798 9650 12850 9662
rect 14926 9714 14978 9726
rect 14926 9650 14978 9662
rect 16830 9714 16882 9726
rect 16830 9650 16882 9662
rect 17838 9714 17890 9726
rect 17838 9650 17890 9662
rect 18398 9714 18450 9726
rect 18398 9650 18450 9662
rect 19518 9714 19570 9726
rect 19518 9650 19570 9662
rect 19630 9714 19682 9726
rect 19630 9650 19682 9662
rect 19854 9714 19906 9726
rect 19854 9650 19906 9662
rect 20302 9714 20354 9726
rect 20302 9650 20354 9662
rect 28814 9714 28866 9726
rect 37550 9714 37602 9726
rect 31154 9662 31166 9714
rect 31218 9662 31230 9714
rect 31490 9662 31502 9714
rect 31554 9662 31566 9714
rect 28814 9650 28866 9662
rect 37550 9650 37602 9662
rect 38782 9714 38834 9726
rect 38782 9650 38834 9662
rect 39006 9714 39058 9726
rect 39006 9650 39058 9662
rect 39566 9714 39618 9726
rect 39566 9650 39618 9662
rect 2942 9602 2994 9614
rect 2942 9538 2994 9550
rect 3950 9602 4002 9614
rect 3950 9538 4002 9550
rect 4174 9602 4226 9614
rect 4174 9538 4226 9550
rect 6526 9602 6578 9614
rect 6526 9538 6578 9550
rect 8430 9602 8482 9614
rect 8430 9538 8482 9550
rect 9998 9602 10050 9614
rect 9998 9538 10050 9550
rect 10894 9602 10946 9614
rect 10894 9538 10946 9550
rect 11118 9602 11170 9614
rect 11118 9538 11170 9550
rect 13022 9602 13074 9614
rect 13022 9538 13074 9550
rect 15038 9602 15090 9614
rect 15038 9538 15090 9550
rect 17054 9602 17106 9614
rect 17054 9538 17106 9550
rect 20526 9602 20578 9614
rect 20526 9538 20578 9550
rect 21758 9602 21810 9614
rect 21758 9538 21810 9550
rect 21982 9602 22034 9614
rect 21982 9538 22034 9550
rect 28590 9602 28642 9614
rect 35870 9602 35922 9614
rect 31826 9550 31838 9602
rect 31890 9550 31902 9602
rect 28590 9538 28642 9550
rect 35870 9538 35922 9550
rect 36094 9602 36146 9614
rect 36094 9538 36146 9550
rect 36654 9602 36706 9614
rect 36654 9538 36706 9550
rect 39678 9602 39730 9614
rect 39678 9538 39730 9550
rect 1344 9434 42560 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 42560 9434
rect 1344 9348 42560 9382
rect 5406 9266 5458 9278
rect 5406 9202 5458 9214
rect 6526 9266 6578 9278
rect 6526 9202 6578 9214
rect 7086 9266 7138 9278
rect 7086 9202 7138 9214
rect 7198 9266 7250 9278
rect 7198 9202 7250 9214
rect 9998 9266 10050 9278
rect 9998 9202 10050 9214
rect 10110 9266 10162 9278
rect 10110 9202 10162 9214
rect 11678 9266 11730 9278
rect 11678 9202 11730 9214
rect 13470 9266 13522 9278
rect 13470 9202 13522 9214
rect 14702 9266 14754 9278
rect 14702 9202 14754 9214
rect 15262 9266 15314 9278
rect 15262 9202 15314 9214
rect 16158 9266 16210 9278
rect 16158 9202 16210 9214
rect 16270 9266 16322 9278
rect 16270 9202 16322 9214
rect 17838 9266 17890 9278
rect 17838 9202 17890 9214
rect 19182 9266 19234 9278
rect 19182 9202 19234 9214
rect 19294 9266 19346 9278
rect 19294 9202 19346 9214
rect 20414 9266 20466 9278
rect 20414 9202 20466 9214
rect 20638 9266 20690 9278
rect 20638 9202 20690 9214
rect 32062 9266 32114 9278
rect 32062 9202 32114 9214
rect 32622 9266 32674 9278
rect 32622 9202 32674 9214
rect 33518 9266 33570 9278
rect 33518 9202 33570 9214
rect 33742 9266 33794 9278
rect 33742 9202 33794 9214
rect 39230 9266 39282 9278
rect 39230 9202 39282 9214
rect 39790 9266 39842 9278
rect 39790 9202 39842 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 41470 9266 41522 9278
rect 41470 9202 41522 9214
rect 41918 9266 41970 9278
rect 41918 9202 41970 9214
rect 6414 9154 6466 9166
rect 3938 9102 3950 9154
rect 4002 9102 4014 9154
rect 6414 9090 6466 9102
rect 7534 9154 7586 9166
rect 7534 9090 7586 9102
rect 8318 9154 8370 9166
rect 8318 9090 8370 9102
rect 8766 9154 8818 9166
rect 8766 9090 8818 9102
rect 11118 9154 11170 9166
rect 11118 9090 11170 9102
rect 12238 9154 12290 9166
rect 12238 9090 12290 9102
rect 13358 9154 13410 9166
rect 16718 9154 16770 9166
rect 14018 9102 14030 9154
rect 14082 9102 14094 9154
rect 13358 9090 13410 9102
rect 16718 9090 16770 9102
rect 18062 9154 18114 9166
rect 18062 9090 18114 9102
rect 18286 9154 18338 9166
rect 18286 9090 18338 9102
rect 29486 9154 29538 9166
rect 29486 9090 29538 9102
rect 30270 9154 30322 9166
rect 30270 9090 30322 9102
rect 31278 9154 31330 9166
rect 38110 9154 38162 9166
rect 35410 9102 35422 9154
rect 35474 9102 35486 9154
rect 31278 9090 31330 9102
rect 38110 9090 38162 9102
rect 5854 9042 5906 9054
rect 4722 8990 4734 9042
rect 4786 8990 4798 9042
rect 5854 8978 5906 8990
rect 6302 9042 6354 9054
rect 6302 8978 6354 8990
rect 7310 9042 7362 9054
rect 9886 9042 9938 9054
rect 15822 9042 15874 9054
rect 17614 9042 17666 9054
rect 21422 9042 21474 9054
rect 33854 9042 33906 9054
rect 38222 9042 38274 9054
rect 8530 8990 8542 9042
rect 8594 8990 8606 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 12674 8990 12686 9042
rect 12738 8990 12750 9042
rect 14242 8990 14254 9042
rect 14306 8990 14318 9042
rect 15474 8990 15486 9042
rect 15538 8990 15550 9042
rect 16482 8990 16494 9042
rect 16546 8990 16558 9042
rect 20850 8990 20862 9042
rect 20914 8990 20926 9042
rect 22082 8990 22094 9042
rect 22146 8990 22158 9042
rect 28578 8990 28590 9042
rect 28642 8990 28654 9042
rect 29250 8990 29262 9042
rect 29314 8990 29326 9042
rect 30930 8990 30942 9042
rect 30994 8990 31006 9042
rect 34738 8990 34750 9042
rect 34802 8990 34814 9042
rect 7310 8978 7362 8990
rect 9886 8978 9938 8990
rect 15822 8978 15874 8990
rect 17614 8978 17666 8990
rect 21422 8978 21474 8990
rect 33854 8978 33906 8990
rect 38222 8978 38274 8990
rect 38446 9042 38498 9054
rect 38658 8990 38670 9042
rect 38722 8990 38734 9042
rect 38446 8978 38498 8990
rect 5294 8930 5346 8942
rect 1810 8878 1822 8930
rect 1874 8878 1886 8930
rect 5294 8866 5346 8878
rect 13582 8930 13634 8942
rect 19854 8930 19906 8942
rect 15362 8878 15374 8930
rect 15426 8878 15438 8930
rect 13582 8866 13634 8878
rect 19854 8866 19906 8878
rect 20750 8930 20802 8942
rect 31838 8930 31890 8942
rect 39342 8930 39394 8942
rect 22754 8878 22766 8930
rect 22818 8878 22830 8930
rect 24882 8878 24894 8930
rect 24946 8878 24958 8930
rect 25666 8878 25678 8930
rect 25730 8878 25742 8930
rect 27794 8878 27806 8930
rect 27858 8878 27870 8930
rect 30258 8878 30270 8930
rect 30322 8878 30334 8930
rect 37538 8878 37550 8930
rect 37602 8878 37614 8930
rect 20750 8866 20802 8878
rect 31838 8866 31890 8878
rect 39342 8866 39394 8878
rect 40686 8930 40738 8942
rect 40686 8866 40738 8878
rect 8206 8818 8258 8830
rect 8206 8754 8258 8766
rect 13806 8818 13858 8830
rect 13806 8754 13858 8766
rect 19406 8818 19458 8830
rect 19406 8754 19458 8766
rect 30046 8818 30098 8830
rect 30046 8754 30098 8766
rect 30942 8818 30994 8830
rect 30942 8754 30994 8766
rect 32174 8818 32226 8830
rect 32386 8766 32398 8818
rect 32450 8815 32462 8818
rect 33058 8815 33070 8818
rect 32450 8769 33070 8815
rect 32450 8766 32462 8769
rect 33058 8766 33070 8769
rect 33122 8766 33134 8818
rect 32174 8754 32226 8766
rect 1344 8650 42560 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 42560 8650
rect 1344 8564 42560 8598
rect 1934 8482 1986 8494
rect 1934 8418 1986 8430
rect 14142 8482 14194 8494
rect 14142 8418 14194 8430
rect 15262 8482 15314 8494
rect 15262 8418 15314 8430
rect 35534 8482 35586 8494
rect 35534 8418 35586 8430
rect 37550 8482 37602 8494
rect 37550 8418 37602 8430
rect 1822 8370 1874 8382
rect 1822 8306 1874 8318
rect 3054 8370 3106 8382
rect 3054 8306 3106 8318
rect 5966 8370 6018 8382
rect 5966 8306 6018 8318
rect 7086 8370 7138 8382
rect 7086 8306 7138 8318
rect 8206 8370 8258 8382
rect 13806 8370 13858 8382
rect 12786 8318 12798 8370
rect 12850 8318 12862 8370
rect 8206 8306 8258 8318
rect 13806 8306 13858 8318
rect 15150 8370 15202 8382
rect 15150 8306 15202 8318
rect 15822 8370 15874 8382
rect 15822 8306 15874 8318
rect 20526 8370 20578 8382
rect 20526 8306 20578 8318
rect 21982 8370 22034 8382
rect 21982 8306 22034 8318
rect 31054 8370 31106 8382
rect 31054 8306 31106 8318
rect 31166 8370 31218 8382
rect 31166 8306 31218 8318
rect 31838 8370 31890 8382
rect 31838 8306 31890 8318
rect 34526 8370 34578 8382
rect 34526 8306 34578 8318
rect 39566 8370 39618 8382
rect 39566 8306 39618 8318
rect 40126 8370 40178 8382
rect 40126 8306 40178 8318
rect 41582 8370 41634 8382
rect 41582 8306 41634 8318
rect 3950 8258 4002 8270
rect 2482 8206 2494 8258
rect 2546 8206 2558 8258
rect 2706 8206 2718 8258
rect 2770 8206 2782 8258
rect 3950 8194 4002 8206
rect 6190 8258 6242 8270
rect 6190 8194 6242 8206
rect 6302 8258 6354 8270
rect 13918 8258 13970 8270
rect 14702 8258 14754 8270
rect 9314 8206 9326 8258
rect 9378 8206 9390 8258
rect 9986 8206 9998 8258
rect 10050 8206 10062 8258
rect 14354 8206 14366 8258
rect 14418 8206 14430 8258
rect 6302 8194 6354 8206
rect 13918 8194 13970 8206
rect 14702 8194 14754 8206
rect 16046 8258 16098 8270
rect 16046 8194 16098 8206
rect 17166 8258 17218 8270
rect 19294 8258 19346 8270
rect 17602 8206 17614 8258
rect 17666 8206 17678 8258
rect 17166 8194 17218 8206
rect 19294 8194 19346 8206
rect 19518 8258 19570 8270
rect 19518 8194 19570 8206
rect 20302 8258 20354 8270
rect 20302 8194 20354 8206
rect 22206 8258 22258 8270
rect 29822 8258 29874 8270
rect 23090 8206 23102 8258
rect 23154 8206 23166 8258
rect 22206 8194 22258 8206
rect 29822 8194 29874 8206
rect 30382 8258 30434 8270
rect 32510 8258 32562 8270
rect 31378 8206 31390 8258
rect 31442 8206 31454 8258
rect 30382 8194 30434 8206
rect 32510 8194 32562 8206
rect 35646 8258 35698 8270
rect 35646 8194 35698 8206
rect 36206 8258 36258 8270
rect 36206 8194 36258 8206
rect 36542 8258 36594 8270
rect 36542 8194 36594 8206
rect 38670 8258 38722 8270
rect 39218 8206 39230 8258
rect 39282 8206 39294 8258
rect 38670 8194 38722 8206
rect 2942 8146 2994 8158
rect 2942 8082 2994 8094
rect 3502 8146 3554 8158
rect 3502 8082 3554 8094
rect 4734 8146 4786 8158
rect 4734 8082 4786 8094
rect 5070 8146 5122 8158
rect 5070 8082 5122 8094
rect 5742 8146 5794 8158
rect 5742 8082 5794 8094
rect 6638 8146 6690 8158
rect 13694 8146 13746 8158
rect 10658 8094 10670 8146
rect 10722 8094 10734 8146
rect 6638 8082 6690 8094
rect 13694 8082 13746 8094
rect 16942 8146 16994 8158
rect 16942 8082 16994 8094
rect 18846 8146 18898 8158
rect 19742 8146 19794 8158
rect 19058 8094 19070 8146
rect 19122 8094 19134 8146
rect 18846 8082 18898 8094
rect 19742 8082 19794 8094
rect 20862 8146 20914 8158
rect 20862 8082 20914 8094
rect 21870 8146 21922 8158
rect 21870 8082 21922 8094
rect 22430 8146 22482 8158
rect 33966 8146 34018 8158
rect 26786 8094 26798 8146
rect 26850 8094 26862 8146
rect 22430 8082 22482 8094
rect 33966 8082 34018 8094
rect 34638 8146 34690 8158
rect 34638 8082 34690 8094
rect 34750 8146 34802 8158
rect 34750 8082 34802 8094
rect 38558 8146 38610 8158
rect 38558 8082 38610 8094
rect 40238 8146 40290 8158
rect 40238 8082 40290 8094
rect 41134 8146 41186 8158
rect 41134 8082 41186 8094
rect 3726 8034 3778 8046
rect 3726 7970 3778 7982
rect 3838 8034 3890 8046
rect 3838 7970 3890 7982
rect 4062 8034 4114 8046
rect 4062 7970 4114 7982
rect 4846 8034 4898 8046
rect 4846 7970 4898 7982
rect 5630 8034 5682 8046
rect 5630 7970 5682 7982
rect 7646 8034 7698 8046
rect 7646 7970 7698 7982
rect 8766 8034 8818 8046
rect 8766 7970 8818 7982
rect 8878 8034 8930 8046
rect 8878 7970 8930 7982
rect 8990 8034 9042 8046
rect 17278 8034 17330 8046
rect 16370 7982 16382 8034
rect 16434 7982 16446 8034
rect 8990 7970 9042 7982
rect 17278 7970 17330 7982
rect 17390 8034 17442 8046
rect 17390 7970 17442 7982
rect 18286 8034 18338 8046
rect 18286 7970 18338 7982
rect 19854 8034 19906 8046
rect 19854 7970 19906 7982
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 28702 8034 28754 8046
rect 28702 7970 28754 7982
rect 30270 8034 30322 8046
rect 30270 7970 30322 7982
rect 30494 8034 30546 8046
rect 30494 7970 30546 7982
rect 32622 8034 32674 8046
rect 32622 7970 32674 7982
rect 32734 8034 32786 8046
rect 32734 7970 32786 7982
rect 32958 8034 33010 8046
rect 32958 7970 33010 7982
rect 33742 8034 33794 8046
rect 33742 7970 33794 7982
rect 33854 8034 33906 8046
rect 33854 7970 33906 7982
rect 35534 8034 35586 8046
rect 35534 7970 35586 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 37662 8034 37714 8046
rect 37662 7970 37714 7982
rect 37774 8034 37826 8046
rect 37774 7970 37826 7982
rect 38334 8034 38386 8046
rect 38334 7970 38386 7982
rect 39454 8034 39506 8046
rect 39454 7970 39506 7982
rect 40686 8034 40738 8046
rect 40686 7970 40738 7982
rect 42030 8034 42082 8046
rect 42030 7970 42082 7982
rect 1344 7866 42560 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 42560 7866
rect 1344 7780 42560 7814
rect 7086 7698 7138 7710
rect 7086 7634 7138 7646
rect 7310 7698 7362 7710
rect 7310 7634 7362 7646
rect 9102 7698 9154 7710
rect 9102 7634 9154 7646
rect 10782 7698 10834 7710
rect 10782 7634 10834 7646
rect 11006 7698 11058 7710
rect 11006 7634 11058 7646
rect 17614 7698 17666 7710
rect 17614 7634 17666 7646
rect 17726 7698 17778 7710
rect 17726 7634 17778 7646
rect 17950 7698 18002 7710
rect 17950 7634 18002 7646
rect 20302 7698 20354 7710
rect 20302 7634 20354 7646
rect 24446 7698 24498 7710
rect 24446 7634 24498 7646
rect 25790 7698 25842 7710
rect 25790 7634 25842 7646
rect 27582 7698 27634 7710
rect 27582 7634 27634 7646
rect 27694 7698 27746 7710
rect 27694 7634 27746 7646
rect 27806 7698 27858 7710
rect 27806 7634 27858 7646
rect 38334 7698 38386 7710
rect 38334 7634 38386 7646
rect 41806 7698 41858 7710
rect 41806 7634 41858 7646
rect 7982 7586 8034 7598
rect 18174 7586 18226 7598
rect 3938 7534 3950 7586
rect 4002 7534 4014 7586
rect 10434 7534 10446 7586
rect 10498 7534 10510 7586
rect 13122 7534 13134 7586
rect 13186 7534 13198 7586
rect 7982 7522 8034 7534
rect 18174 7522 18226 7534
rect 25902 7586 25954 7598
rect 31950 7586 32002 7598
rect 29138 7534 29150 7586
rect 29202 7534 29214 7586
rect 25902 7522 25954 7534
rect 31950 7522 32002 7534
rect 32286 7586 32338 7598
rect 32286 7522 32338 7534
rect 32510 7586 32562 7598
rect 32510 7522 32562 7534
rect 33630 7586 33682 7598
rect 33630 7522 33682 7534
rect 33854 7586 33906 7598
rect 38222 7586 38274 7598
rect 35522 7534 35534 7586
rect 35586 7534 35598 7586
rect 33854 7522 33906 7534
rect 38222 7522 38274 7534
rect 5518 7474 5570 7486
rect 6862 7474 6914 7486
rect 4722 7422 4734 7474
rect 4786 7422 4798 7474
rect 6178 7422 6190 7474
rect 6242 7422 6254 7474
rect 5518 7410 5570 7422
rect 6862 7410 6914 7422
rect 6974 7474 7026 7486
rect 6974 7410 7026 7422
rect 8206 7474 8258 7486
rect 8206 7410 8258 7422
rect 8430 7474 8482 7486
rect 19070 7474 19122 7486
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 16594 7422 16606 7474
rect 16658 7422 16670 7474
rect 18722 7422 18734 7474
rect 18786 7422 18798 7474
rect 8430 7410 8482 7422
rect 19070 7410 19122 7422
rect 19630 7474 19682 7486
rect 27134 7474 27186 7486
rect 20850 7422 20862 7474
rect 20914 7422 20926 7474
rect 24210 7422 24222 7474
rect 24274 7422 24286 7474
rect 28466 7422 28478 7474
rect 28530 7422 28542 7474
rect 34738 7422 34750 7474
rect 34802 7422 34814 7474
rect 40114 7422 40126 7474
rect 40178 7422 40190 7474
rect 19630 7410 19682 7422
rect 27134 7410 27186 7422
rect 5966 7362 6018 7374
rect 1810 7310 1822 7362
rect 1874 7310 1886 7362
rect 5966 7298 6018 7310
rect 9774 7362 9826 7374
rect 19406 7362 19458 7374
rect 10658 7310 10670 7362
rect 10722 7310 10734 7362
rect 9774 7298 9826 7310
rect 19406 7298 19458 7310
rect 19518 7362 19570 7374
rect 26686 7362 26738 7374
rect 32062 7362 32114 7374
rect 40686 7362 40738 7374
rect 21522 7310 21534 7362
rect 21586 7310 21598 7362
rect 23650 7310 23662 7362
rect 23714 7310 23726 7362
rect 31266 7310 31278 7362
rect 31330 7310 31342 7362
rect 33954 7310 33966 7362
rect 34018 7310 34030 7362
rect 37650 7310 37662 7362
rect 37714 7310 37726 7362
rect 39218 7310 39230 7362
rect 39282 7310 39294 7362
rect 19518 7298 19570 7310
rect 26686 7298 26738 7310
rect 32062 7298 32114 7310
rect 40686 7298 40738 7310
rect 41694 7362 41746 7374
rect 41694 7298 41746 7310
rect 5406 7250 5458 7262
rect 5406 7186 5458 7198
rect 5742 7250 5794 7262
rect 5742 7186 5794 7198
rect 8654 7250 8706 7262
rect 8654 7186 8706 7198
rect 19182 7250 19234 7262
rect 19182 7186 19234 7198
rect 24558 7250 24610 7262
rect 24558 7186 24610 7198
rect 25678 7250 25730 7262
rect 25678 7186 25730 7198
rect 26574 7250 26626 7262
rect 26574 7186 26626 7198
rect 40798 7250 40850 7262
rect 40798 7186 40850 7198
rect 41582 7250 41634 7262
rect 41582 7186 41634 7198
rect 1344 7082 42560 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 42560 7082
rect 1344 6996 42560 7030
rect 15598 6914 15650 6926
rect 15598 6850 15650 6862
rect 17054 6914 17106 6926
rect 29598 6914 29650 6926
rect 28690 6862 28702 6914
rect 28754 6911 28766 6914
rect 28914 6911 28926 6914
rect 28754 6865 28926 6911
rect 28754 6862 28766 6865
rect 28914 6862 28926 6865
rect 28978 6862 28990 6914
rect 17054 6850 17106 6862
rect 29598 6850 29650 6862
rect 29934 6914 29986 6926
rect 29934 6850 29986 6862
rect 36318 6914 36370 6926
rect 36318 6850 36370 6862
rect 5966 6802 6018 6814
rect 4162 6750 4174 6802
rect 4226 6750 4238 6802
rect 5966 6738 6018 6750
rect 7422 6802 7474 6814
rect 15262 6802 15314 6814
rect 11554 6750 11566 6802
rect 11618 6750 11630 6802
rect 7422 6738 7474 6750
rect 15262 6738 15314 6750
rect 20526 6802 20578 6814
rect 36766 6802 36818 6814
rect 23538 6750 23550 6802
rect 23602 6750 23614 6802
rect 31938 6750 31950 6802
rect 32002 6750 32014 6802
rect 34066 6750 34078 6802
rect 34130 6750 34142 6802
rect 36082 6750 36094 6802
rect 36146 6750 36158 6802
rect 20526 6738 20578 6750
rect 36766 6738 36818 6750
rect 37774 6802 37826 6814
rect 37774 6738 37826 6750
rect 41246 6802 41298 6814
rect 41246 6738 41298 6750
rect 4734 6690 4786 6702
rect 4734 6626 4786 6638
rect 6190 6690 6242 6702
rect 7534 6690 7586 6702
rect 6402 6638 6414 6690
rect 6466 6638 6478 6690
rect 6626 6638 6638 6690
rect 6690 6638 6702 6690
rect 6190 6626 6242 6638
rect 7534 6626 7586 6638
rect 9550 6690 9602 6702
rect 10334 6690 10386 6702
rect 9986 6638 9998 6690
rect 10050 6638 10062 6690
rect 9550 6626 9602 6638
rect 10334 6626 10386 6638
rect 10446 6690 10498 6702
rect 10446 6626 10498 6638
rect 10558 6690 10610 6702
rect 12686 6690 12738 6702
rect 15150 6690 15202 6702
rect 12226 6638 12238 6690
rect 12290 6638 12302 6690
rect 14354 6638 14366 6690
rect 14418 6638 14430 6690
rect 10558 6626 10610 6638
rect 12686 6626 12738 6638
rect 15150 6626 15202 6638
rect 15374 6690 15426 6702
rect 15374 6626 15426 6638
rect 15710 6690 15762 6702
rect 15710 6626 15762 6638
rect 16494 6690 16546 6702
rect 16494 6626 16546 6638
rect 17278 6690 17330 6702
rect 17278 6626 17330 6638
rect 18622 6690 18674 6702
rect 18622 6626 18674 6638
rect 18846 6690 18898 6702
rect 20414 6690 20466 6702
rect 20178 6638 20190 6690
rect 20242 6638 20254 6690
rect 18846 6626 18898 6638
rect 20414 6626 20466 6638
rect 20750 6690 20802 6702
rect 20750 6626 20802 6638
rect 22318 6690 22370 6702
rect 30606 6690 30658 6702
rect 34862 6690 34914 6702
rect 28242 6638 28254 6690
rect 28306 6638 28318 6690
rect 31154 6638 31166 6690
rect 31218 6638 31230 6690
rect 22318 6626 22370 6638
rect 30606 6626 30658 6638
rect 34862 6626 34914 6638
rect 35086 6690 35138 6702
rect 35086 6626 35138 6638
rect 35534 6690 35586 6702
rect 37886 6690 37938 6702
rect 41918 6690 41970 6702
rect 35970 6638 35982 6690
rect 36034 6638 36046 6690
rect 40114 6638 40126 6690
rect 40178 6638 40190 6690
rect 40786 6638 40798 6690
rect 40850 6638 40862 6690
rect 35534 6626 35586 6638
rect 37886 6626 37938 6638
rect 41918 6626 41970 6638
rect 2158 6578 2210 6590
rect 5742 6578 5794 6590
rect 9214 6578 9266 6590
rect 2818 6526 2830 6578
rect 2882 6526 2894 6578
rect 7858 6526 7870 6578
rect 7922 6526 7934 6578
rect 8418 6526 8430 6578
rect 8482 6526 8494 6578
rect 2158 6514 2210 6526
rect 5742 6514 5794 6526
rect 9214 6514 9266 6526
rect 9326 6578 9378 6590
rect 9326 6514 9378 6526
rect 12462 6578 12514 6590
rect 16046 6578 16098 6590
rect 17502 6578 17554 6590
rect 13794 6526 13806 6578
rect 13858 6526 13870 6578
rect 14130 6526 14142 6578
rect 14194 6526 14206 6578
rect 16818 6526 16830 6578
rect 16882 6526 16894 6578
rect 12462 6514 12514 6526
rect 16046 6514 16098 6526
rect 17502 6514 17554 6526
rect 18398 6578 18450 6590
rect 19294 6578 19346 6590
rect 19058 6526 19070 6578
rect 19122 6526 19134 6578
rect 18398 6514 18450 6526
rect 19294 6514 19346 6526
rect 30494 6578 30546 6590
rect 30494 6514 30546 6526
rect 38110 6578 38162 6590
rect 38994 6526 39006 6578
rect 39058 6526 39070 6578
rect 38110 6514 38162 6526
rect 2046 6466 2098 6478
rect 2046 6402 2098 6414
rect 4846 6466 4898 6478
rect 4846 6402 4898 6414
rect 5070 6466 5122 6478
rect 5070 6402 5122 6414
rect 5630 6466 5682 6478
rect 5630 6402 5682 6414
rect 11118 6466 11170 6478
rect 11118 6402 11170 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 12798 6466 12850 6478
rect 18286 6466 18338 6478
rect 16930 6414 16942 6466
rect 16994 6414 17006 6466
rect 12798 6402 12850 6414
rect 18286 6402 18338 6414
rect 20638 6466 20690 6478
rect 20638 6402 20690 6414
rect 21646 6466 21698 6478
rect 21646 6402 21698 6414
rect 21758 6466 21810 6478
rect 21758 6402 21810 6414
rect 21870 6466 21922 6478
rect 21870 6402 21922 6414
rect 28702 6466 28754 6478
rect 28702 6402 28754 6414
rect 29822 6466 29874 6478
rect 29822 6402 29874 6414
rect 35310 6466 35362 6478
rect 35310 6402 35362 6414
rect 37662 6466 37714 6478
rect 37662 6402 37714 6414
rect 42030 6466 42082 6478
rect 42030 6402 42082 6414
rect 1344 6298 42560 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 42560 6298
rect 1344 6212 42560 6246
rect 10334 6130 10386 6142
rect 10334 6066 10386 6078
rect 16942 6130 16994 6142
rect 16942 6066 16994 6078
rect 23774 6130 23826 6142
rect 23774 6066 23826 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 24782 6130 24834 6142
rect 28478 6130 28530 6142
rect 26786 6078 26798 6130
rect 26850 6078 26862 6130
rect 24782 6066 24834 6078
rect 28478 6066 28530 6078
rect 29374 6130 29426 6142
rect 29374 6066 29426 6078
rect 29598 6130 29650 6142
rect 29598 6066 29650 6078
rect 33854 6130 33906 6142
rect 33854 6066 33906 6078
rect 34190 6130 34242 6142
rect 34190 6066 34242 6078
rect 38222 6130 38274 6142
rect 38222 6066 38274 6078
rect 40238 6130 40290 6142
rect 40238 6066 40290 6078
rect 41694 6130 41746 6142
rect 41694 6066 41746 6078
rect 41806 6130 41858 6142
rect 41806 6066 41858 6078
rect 11566 6018 11618 6030
rect 16830 6018 16882 6030
rect 28590 6018 28642 6030
rect 5506 5966 5518 6018
rect 5570 5966 5582 6018
rect 8866 5966 8878 6018
rect 8930 5966 8942 6018
rect 12338 5966 12350 6018
rect 12402 5966 12414 6018
rect 15810 5966 15822 6018
rect 15874 5966 15886 6018
rect 19618 5966 19630 6018
rect 19682 5966 19694 6018
rect 22418 5966 22430 6018
rect 22482 5966 22494 6018
rect 11566 5954 11618 5966
rect 16830 5954 16882 5966
rect 28590 5954 28642 5966
rect 29934 6018 29986 6030
rect 29934 5954 29986 5966
rect 31502 6018 31554 6030
rect 31502 5954 31554 5966
rect 31838 6018 31890 6030
rect 31838 5954 31890 5966
rect 32734 6018 32786 6030
rect 32734 5954 32786 5966
rect 32846 6018 32898 6030
rect 32846 5954 32898 5966
rect 33630 6018 33682 6030
rect 33630 5954 33682 5966
rect 34078 6018 34130 6030
rect 40126 6018 40178 6030
rect 35410 5966 35422 6018
rect 35474 5966 35486 6018
rect 34078 5954 34130 5966
rect 38558 5962 38610 5974
rect 39554 5966 39566 6018
rect 39618 5966 39630 6018
rect 9886 5906 9938 5918
rect 1922 5854 1934 5906
rect 1986 5854 1998 5906
rect 9886 5842 9938 5854
rect 9998 5906 10050 5918
rect 9998 5842 10050 5854
rect 10222 5906 10274 5918
rect 10222 5842 10274 5854
rect 11006 5906 11058 5918
rect 11006 5842 11058 5854
rect 17726 5906 17778 5918
rect 24670 5906 24722 5918
rect 23202 5854 23214 5906
rect 23266 5854 23278 5906
rect 24210 5854 24222 5906
rect 24274 5854 24286 5906
rect 17726 5842 17778 5854
rect 24670 5842 24722 5854
rect 25678 5906 25730 5918
rect 25678 5842 25730 5854
rect 26238 5906 26290 5918
rect 26238 5842 26290 5854
rect 26462 5906 26514 5918
rect 26462 5842 26514 5854
rect 27470 5906 27522 5918
rect 27470 5842 27522 5854
rect 27694 5906 27746 5918
rect 27694 5842 27746 5854
rect 28030 5906 28082 5918
rect 28030 5842 28082 5854
rect 29262 5906 29314 5918
rect 29262 5842 29314 5854
rect 29822 5906 29874 5918
rect 29822 5842 29874 5854
rect 30382 5906 30434 5918
rect 30382 5842 30434 5854
rect 30494 5906 30546 5918
rect 30494 5842 30546 5854
rect 30718 5906 30770 5918
rect 32062 5906 32114 5918
rect 30930 5854 30942 5906
rect 30994 5854 31006 5906
rect 30718 5842 30770 5854
rect 32062 5842 32114 5854
rect 32510 5906 32562 5918
rect 38110 5906 38162 5918
rect 34626 5854 34638 5906
rect 34690 5854 34702 5906
rect 40126 5954 40178 5966
rect 41582 6018 41634 6030
rect 41582 5954 41634 5966
rect 38558 5898 38610 5910
rect 39330 5854 39342 5906
rect 39394 5854 39406 5906
rect 40450 5854 40462 5906
rect 40514 5854 40526 5906
rect 32510 5842 32562 5854
rect 38110 5842 38162 5854
rect 10110 5794 10162 5806
rect 14142 5794 14194 5806
rect 24558 5794 24610 5806
rect 2594 5742 2606 5794
rect 2658 5742 2670 5794
rect 4722 5742 4734 5794
rect 4786 5742 4798 5794
rect 6738 5742 6750 5794
rect 6802 5742 6814 5794
rect 7634 5742 7646 5794
rect 7698 5742 7710 5794
rect 13458 5742 13470 5794
rect 13522 5742 13534 5794
rect 14802 5742 14814 5794
rect 14866 5742 14878 5794
rect 18498 5742 18510 5794
rect 18562 5742 18574 5794
rect 20290 5742 20302 5794
rect 20354 5742 20366 5794
rect 10110 5730 10162 5742
rect 14142 5730 14194 5742
rect 24558 5730 24610 5742
rect 27806 5794 27858 5806
rect 27806 5730 27858 5742
rect 31614 5794 31666 5806
rect 37538 5742 37550 5794
rect 37602 5742 37614 5794
rect 31614 5730 31666 5742
rect 14254 5682 14306 5694
rect 14254 5618 14306 5630
rect 1344 5514 42560 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 42560 5514
rect 1344 5428 42560 5462
rect 5854 5346 5906 5358
rect 5854 5282 5906 5294
rect 12014 5346 12066 5358
rect 33630 5346 33682 5358
rect 20290 5294 20302 5346
rect 20354 5294 20366 5346
rect 12014 5282 12066 5294
rect 33630 5282 33682 5294
rect 35982 5346 36034 5358
rect 35982 5282 36034 5294
rect 36318 5346 36370 5358
rect 36318 5282 36370 5294
rect 1822 5234 1874 5246
rect 1822 5170 1874 5182
rect 2606 5234 2658 5246
rect 14254 5234 14306 5246
rect 33406 5234 33458 5246
rect 36766 5234 36818 5246
rect 37886 5234 37938 5246
rect 4946 5182 4958 5234
rect 5010 5182 5022 5234
rect 6402 5182 6414 5234
rect 6466 5182 6478 5234
rect 8418 5182 8430 5234
rect 8482 5182 8494 5234
rect 10546 5182 10558 5234
rect 10610 5182 10622 5234
rect 14802 5182 14814 5234
rect 14866 5182 14878 5234
rect 17602 5182 17614 5234
rect 17666 5182 17678 5234
rect 19730 5182 19742 5234
rect 19794 5182 19806 5234
rect 24658 5182 24670 5234
rect 24722 5182 24734 5234
rect 26786 5182 26798 5234
rect 26850 5182 26862 5234
rect 30706 5182 30718 5234
rect 30770 5182 30782 5234
rect 32834 5182 32846 5234
rect 32898 5182 32910 5234
rect 33954 5182 33966 5234
rect 34018 5182 34030 5234
rect 37538 5182 37550 5234
rect 37602 5182 37614 5234
rect 2606 5170 2658 5182
rect 14254 5170 14306 5182
rect 33406 5170 33458 5182
rect 36766 5170 36818 5182
rect 37886 5170 37938 5182
rect 38334 5234 38386 5246
rect 41346 5182 41358 5234
rect 41410 5182 41422 5234
rect 38334 5170 38386 5182
rect 12574 5122 12626 5134
rect 23438 5122 23490 5134
rect 34974 5122 35026 5134
rect 2258 5070 2270 5122
rect 2322 5070 2334 5122
rect 11218 5070 11230 5122
rect 11282 5070 11294 5122
rect 16818 5070 16830 5122
rect 16882 5070 16894 5122
rect 20514 5070 20526 5122
rect 20578 5070 20590 5122
rect 23986 5070 23998 5122
rect 24050 5070 24062 5122
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 29922 5070 29934 5122
rect 29986 5070 29998 5122
rect 39890 5070 39902 5122
rect 39954 5070 39966 5122
rect 40674 5070 40686 5122
rect 40738 5070 40750 5122
rect 12574 5058 12626 5070
rect 23438 5058 23490 5070
rect 34974 5058 35026 5070
rect 2494 5010 2546 5022
rect 2494 4946 2546 4958
rect 2718 5010 2770 5022
rect 5742 5010 5794 5022
rect 11902 5010 11954 5022
rect 3826 4958 3838 5010
rect 3890 4958 3902 5010
rect 7410 4958 7422 5010
rect 7474 4958 7486 5010
rect 2718 4946 2770 4958
rect 5742 4946 5794 4958
rect 11902 4946 11954 4958
rect 12126 5010 12178 5022
rect 12126 4946 12178 4958
rect 12350 5010 12402 5022
rect 21870 5010 21922 5022
rect 15922 4958 15934 5010
rect 15986 4958 15998 5010
rect 12350 4946 12402 4958
rect 21870 4946 21922 4958
rect 22430 5010 22482 5022
rect 22430 4946 22482 4958
rect 23102 5010 23154 5022
rect 35086 5010 35138 5022
rect 27458 4958 27470 5010
rect 27522 4958 27534 5010
rect 23102 4946 23154 4958
rect 35086 4946 35138 4958
rect 35422 5010 35474 5022
rect 35422 4946 35474 4958
rect 36094 5010 36146 5022
rect 38994 4958 39006 5010
rect 39058 4958 39070 5010
rect 36094 4946 36146 4958
rect 2830 4898 2882 4910
rect 2830 4834 2882 4846
rect 13694 4898 13746 4910
rect 13694 4834 13746 4846
rect 22094 4898 22146 4910
rect 22094 4834 22146 4846
rect 22206 4898 22258 4910
rect 22206 4834 22258 4846
rect 22318 4898 22370 4910
rect 22318 4834 22370 4846
rect 23214 4898 23266 4910
rect 23214 4834 23266 4846
rect 35310 4898 35362 4910
rect 35310 4834 35362 4846
rect 1344 4730 42560 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 42560 4730
rect 1344 4644 42560 4678
rect 6750 4562 6802 4574
rect 6750 4498 6802 4510
rect 6974 4562 7026 4574
rect 6974 4498 7026 4510
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 29038 4562 29090 4574
rect 29038 4498 29090 4510
rect 32734 4562 32786 4574
rect 32734 4498 32786 4510
rect 40014 4562 40066 4574
rect 40014 4498 40066 4510
rect 40686 4562 40738 4574
rect 40686 4498 40738 4510
rect 6526 4450 6578 4462
rect 9886 4450 9938 4462
rect 1810 4398 1822 4450
rect 1874 4398 1886 4450
rect 7634 4398 7646 4450
rect 7698 4398 7710 4450
rect 6526 4386 6578 4398
rect 9886 4386 9938 4398
rect 18062 4450 18114 4462
rect 24782 4450 24834 4462
rect 32846 4450 32898 4462
rect 21634 4398 21646 4450
rect 21698 4398 21710 4450
rect 26450 4398 26462 4450
rect 26514 4398 26526 4450
rect 18062 4386 18114 4398
rect 24782 4386 24834 4398
rect 32846 4386 32898 4398
rect 33630 4450 33682 4462
rect 40238 4450 40290 4462
rect 35410 4398 35422 4450
rect 35474 4398 35486 4450
rect 33630 4386 33682 4398
rect 40238 4386 40290 4398
rect 41582 4450 41634 4462
rect 41582 4386 41634 4398
rect 18174 4338 18226 4350
rect 2034 4286 2046 4338
rect 2098 4286 2110 4338
rect 5954 4286 5966 4338
rect 6018 4286 6030 4338
rect 10546 4286 10558 4338
rect 10610 4286 10622 4338
rect 13906 4286 13918 4338
rect 13970 4286 13982 4338
rect 14690 4286 14702 4338
rect 14754 4286 14766 4338
rect 18174 4274 18226 4286
rect 18398 4338 18450 4350
rect 18398 4274 18450 4286
rect 18622 4338 18674 4350
rect 31390 4338 31442 4350
rect 22418 4286 22430 4338
rect 22482 4286 22494 4338
rect 23986 4286 23998 4338
rect 24050 4286 24062 4338
rect 25778 4286 25790 4338
rect 25842 4286 25854 4338
rect 30818 4286 30830 4338
rect 30882 4286 30894 4338
rect 18622 4274 18674 4286
rect 31390 4274 31442 4286
rect 31614 4338 31666 4350
rect 31938 4286 31950 4338
rect 32002 4286 32014 4338
rect 32498 4286 32510 4338
rect 32562 4286 32574 4338
rect 33842 4286 33854 4338
rect 33906 4286 33918 4338
rect 34626 4286 34638 4338
rect 34690 4286 34702 4338
rect 39330 4286 39342 4338
rect 39394 4286 39406 4338
rect 41794 4286 41806 4338
rect 41858 4286 41870 4338
rect 31614 4274 31666 4286
rect 3042 4174 3054 4226
rect 3106 4174 3118 4226
rect 5170 4174 5182 4226
rect 5234 4174 5246 4226
rect 8978 4174 8990 4226
rect 9042 4174 9054 4226
rect 11218 4174 11230 4226
rect 11282 4174 11294 4226
rect 13346 4174 13358 4226
rect 13410 4174 13422 4226
rect 16818 4174 16830 4226
rect 16882 4174 16894 4226
rect 19506 4174 19518 4226
rect 19570 4174 19582 4226
rect 23090 4174 23102 4226
rect 23154 4174 23166 4226
rect 28578 4174 28590 4226
rect 28642 4174 28654 4226
rect 29698 4174 29710 4226
rect 29762 4174 29774 4226
rect 37538 4174 37550 4226
rect 37602 4174 37614 4226
rect 38210 4174 38222 4226
rect 38274 4174 38286 4226
rect 7086 4114 7138 4126
rect 7086 4050 7138 4062
rect 18734 4114 18786 4126
rect 18734 4050 18786 4062
rect 24894 4114 24946 4126
rect 24894 4050 24946 4062
rect 39902 4114 39954 4126
rect 39902 4050 39954 4062
rect 1344 3946 42560 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 42560 3946
rect 1344 3860 42560 3894
rect 4958 3778 5010 3790
rect 4958 3714 5010 3726
rect 6862 3778 6914 3790
rect 6862 3714 6914 3726
rect 10110 3778 10162 3790
rect 10110 3714 10162 3726
rect 10334 3778 10386 3790
rect 10334 3714 10386 3726
rect 10558 3778 10610 3790
rect 10558 3714 10610 3726
rect 10670 3778 10722 3790
rect 10670 3714 10722 3726
rect 14030 3778 14082 3790
rect 14030 3714 14082 3726
rect 14254 3778 14306 3790
rect 14254 3714 14306 3726
rect 14478 3778 14530 3790
rect 14478 3714 14530 3726
rect 17726 3778 17778 3790
rect 17726 3714 17778 3726
rect 23550 3778 23602 3790
rect 23550 3714 23602 3726
rect 23886 3778 23938 3790
rect 23886 3714 23938 3726
rect 41918 3778 41970 3790
rect 41918 3714 41970 3726
rect 4846 3666 4898 3678
rect 6750 3666 6802 3678
rect 14590 3666 14642 3678
rect 24446 3666 24498 3678
rect 40910 3666 40962 3678
rect 4162 3614 4174 3666
rect 4226 3614 4238 3666
rect 5842 3614 5854 3666
rect 5906 3614 5918 3666
rect 8866 3614 8878 3666
rect 8930 3614 8942 3666
rect 12786 3614 12798 3666
rect 12850 3614 12862 3666
rect 15474 3614 15486 3666
rect 15538 3614 15550 3666
rect 19170 3614 19182 3666
rect 19234 3614 19246 3666
rect 21522 3614 21534 3666
rect 21586 3614 21598 3666
rect 27794 3614 27806 3666
rect 27858 3614 27870 3666
rect 29922 3614 29934 3666
rect 29986 3614 29998 3666
rect 33842 3614 33854 3666
rect 33906 3614 33918 3666
rect 35634 3614 35646 3666
rect 35698 3614 35710 3666
rect 41570 3614 41582 3666
rect 41634 3614 41646 3666
rect 4846 3602 4898 3614
rect 6750 3602 6802 3614
rect 14590 3602 14642 3614
rect 24446 3602 24498 3614
rect 40910 3602 40962 3614
rect 5966 3554 6018 3566
rect 17614 3554 17666 3566
rect 6178 3502 6190 3554
rect 6242 3502 6254 3554
rect 5966 3490 6018 3502
rect 17614 3490 17666 3502
rect 18286 3554 18338 3566
rect 18286 3490 18338 3502
rect 18622 3554 18674 3566
rect 26338 3502 26350 3554
rect 26402 3502 26414 3554
rect 27234 3502 27246 3554
rect 27298 3502 27310 3554
rect 29474 3502 29486 3554
rect 29538 3502 29550 3554
rect 32274 3502 32286 3554
rect 32338 3502 32350 3554
rect 33170 3502 33182 3554
rect 33234 3502 33246 3554
rect 34962 3502 34974 3554
rect 35026 3502 35038 3554
rect 38322 3502 38334 3554
rect 38386 3502 38398 3554
rect 40114 3502 40126 3554
rect 40178 3502 40190 3554
rect 18622 3490 18674 3502
rect 13918 3442 13970 3454
rect 23774 3442 23826 3454
rect 41694 3442 41746 3454
rect 2258 3390 2270 3442
rect 2322 3390 2334 3442
rect 7858 3390 7870 3442
rect 7922 3390 7934 3442
rect 11666 3390 11678 3442
rect 11730 3390 11742 3442
rect 16594 3390 16606 3442
rect 16658 3390 16670 3442
rect 20178 3390 20190 3442
rect 20242 3390 20254 3442
rect 22530 3390 22542 3442
rect 22594 3390 22606 3442
rect 25442 3390 25454 3442
rect 25506 3390 25518 3442
rect 31154 3390 31166 3442
rect 31218 3390 31230 3442
rect 37202 3390 37214 3442
rect 37266 3390 37278 3442
rect 38994 3390 39006 3442
rect 39058 3390 39070 3442
rect 13918 3378 13970 3390
rect 23774 3378 23826 3390
rect 41694 3378 41746 3390
rect 6414 3330 6466 3342
rect 6414 3266 6466 3278
rect 10222 3330 10274 3342
rect 10222 3266 10274 3278
rect 17726 3330 17778 3342
rect 17726 3266 17778 3278
rect 18510 3330 18562 3342
rect 18510 3266 18562 3278
rect 1344 3162 42560 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 42560 3162
rect 1344 3076 42560 3110
<< via1 >>
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 2494 25454 2546 25506
rect 2942 25230 2994 25282
rect 5070 25230 5122 25282
rect 5742 25230 5794 25282
rect 6190 25230 6242 25282
rect 6974 25230 7026 25282
rect 7422 25230 7474 25282
rect 7870 25230 7922 25282
rect 9550 25230 9602 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2270 24670 2322 24722
rect 6862 24670 6914 24722
rect 1822 24558 1874 24610
rect 2718 24558 2770 24610
rect 3278 24558 3330 24610
rect 4062 24558 4114 24610
rect 4510 24558 4562 24610
rect 5070 24558 5122 24610
rect 5518 24558 5570 24610
rect 5966 24558 6018 24610
rect 6414 24558 6466 24610
rect 7310 24558 7362 24610
rect 7646 24558 7698 24610
rect 8206 24558 8258 24610
rect 8654 24558 8706 24610
rect 9102 24558 9154 24610
rect 9998 24558 10050 24610
rect 10670 24558 10722 24610
rect 11118 24558 11170 24610
rect 8094 24446 8146 24498
rect 9102 24446 9154 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 8766 24110 8818 24162
rect 9550 24110 9602 24162
rect 8654 23998 8706 24050
rect 9102 23998 9154 24050
rect 11230 23998 11282 24050
rect 12238 23998 12290 24050
rect 14030 23998 14082 24050
rect 14478 23998 14530 24050
rect 15038 23998 15090 24050
rect 13582 23886 13634 23938
rect 3726 23774 3778 23826
rect 5742 23774 5794 23826
rect 8318 23774 8370 23826
rect 1934 23662 1986 23714
rect 2382 23662 2434 23714
rect 2830 23662 2882 23714
rect 3278 23662 3330 23714
rect 4174 23662 4226 23714
rect 4622 23662 4674 23714
rect 4958 23662 5010 23714
rect 6302 23662 6354 23714
rect 6862 23662 6914 23714
rect 7422 23662 7474 23714
rect 7758 23662 7810 23714
rect 9662 23662 9714 23714
rect 10110 23662 10162 23714
rect 10894 23662 10946 23714
rect 11902 23662 11954 23714
rect 12686 23662 12738 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 2158 23326 2210 23378
rect 10222 23102 10274 23154
rect 13022 23102 13074 23154
rect 16830 23102 16882 23154
rect 1822 22990 1874 23042
rect 2606 22990 2658 23042
rect 3166 22990 3218 23042
rect 3614 22990 3666 23042
rect 3950 22990 4002 23042
rect 4398 22990 4450 23042
rect 4846 22990 4898 23042
rect 5518 22990 5570 23042
rect 6190 22990 6242 23042
rect 6526 22990 6578 23042
rect 7086 22990 7138 23042
rect 7422 22990 7474 23042
rect 7870 22990 7922 23042
rect 8542 22990 8594 23042
rect 9102 22990 9154 23042
rect 9662 22990 9714 23042
rect 10670 22990 10722 23042
rect 11342 22990 11394 23042
rect 12014 22990 12066 23042
rect 12462 22990 12514 23042
rect 13470 22990 13522 23042
rect 13806 22990 13858 23042
rect 14702 22990 14754 23042
rect 15150 22990 15202 23042
rect 15486 22990 15538 23042
rect 16046 22990 16098 23042
rect 16494 22990 16546 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3950 22542 4002 22594
rect 4958 22542 5010 22594
rect 1822 22430 1874 22482
rect 2718 22430 2770 22482
rect 3054 22430 3106 22482
rect 4398 22430 4450 22482
rect 4846 22430 4898 22482
rect 11342 22430 11394 22482
rect 17390 22430 17442 22482
rect 17838 22430 17890 22482
rect 39118 22318 39170 22370
rect 10110 22206 10162 22258
rect 16494 22206 16546 22258
rect 40014 22206 40066 22258
rect 2158 22094 2210 22146
rect 3614 22094 3666 22146
rect 4062 22094 4114 22146
rect 6078 22094 6130 22146
rect 6414 22094 6466 22146
rect 6862 22094 6914 22146
rect 7758 22094 7810 22146
rect 8094 22094 8146 22146
rect 8542 22094 8594 22146
rect 8990 22094 9042 22146
rect 9550 22094 9602 22146
rect 10446 22094 10498 22146
rect 11006 22094 11058 22146
rect 11790 22094 11842 22146
rect 12350 22094 12402 22146
rect 12910 22094 12962 22146
rect 13694 22094 13746 22146
rect 14142 22094 14194 22146
rect 14926 22094 14978 22146
rect 15374 22094 15426 22146
rect 16158 22094 16210 22146
rect 16942 22094 16994 22146
rect 18286 22094 18338 22146
rect 40574 22094 40626 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2942 21758 2994 21810
rect 4734 21758 4786 21810
rect 5742 21758 5794 21810
rect 6190 21758 6242 21810
rect 7982 21758 8034 21810
rect 10110 21758 10162 21810
rect 10558 21758 10610 21810
rect 11006 21758 11058 21810
rect 14030 21758 14082 21810
rect 16942 21758 16994 21810
rect 17614 21758 17666 21810
rect 19406 21758 19458 21810
rect 4286 21646 4338 21698
rect 16046 21646 16098 21698
rect 16494 21646 16546 21698
rect 3838 21534 3890 21586
rect 5406 21534 5458 21586
rect 2158 21422 2210 21474
rect 2606 21422 2658 21474
rect 3502 21422 3554 21474
rect 6750 21422 6802 21474
rect 7086 21422 7138 21474
rect 7534 21422 7586 21474
rect 8542 21422 8594 21474
rect 9102 21422 9154 21474
rect 9662 21422 9714 21474
rect 11454 21422 11506 21474
rect 12014 21422 12066 21474
rect 12350 21422 12402 21474
rect 13246 21422 13298 21474
rect 13694 21422 13746 21474
rect 14478 21422 14530 21474
rect 14926 21422 14978 21474
rect 15598 21422 15650 21474
rect 18174 21422 18226 21474
rect 18510 21422 18562 21474
rect 18958 21422 19010 21474
rect 2830 21310 2882 21362
rect 3614 21310 3666 21362
rect 8542 21310 8594 21362
rect 8878 21310 8930 21362
rect 9662 21310 9714 21362
rect 10782 21310 10834 21362
rect 11454 21310 11506 21362
rect 12350 21310 12402 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 1934 20974 1986 21026
rect 2494 20974 2546 21026
rect 13806 20974 13858 21026
rect 14590 20974 14642 21026
rect 2382 20862 2434 20914
rect 5630 20862 5682 20914
rect 7086 20862 7138 20914
rect 8990 20862 9042 20914
rect 11902 20862 11954 20914
rect 2046 20638 2098 20690
rect 7982 20638 8034 20690
rect 19630 20638 19682 20690
rect 2830 20526 2882 20578
rect 3502 20526 3554 20578
rect 3950 20526 4002 20578
rect 4622 20526 4674 20578
rect 5070 20526 5122 20578
rect 6302 20526 6354 20578
rect 6638 20526 6690 20578
rect 7646 20526 7698 20578
rect 8542 20526 8594 20578
rect 9438 20526 9490 20578
rect 10222 20526 10274 20578
rect 10670 20526 10722 20578
rect 11454 20526 11506 20578
rect 12462 20526 12514 20578
rect 12910 20526 12962 20578
rect 13582 20526 13634 20578
rect 14142 20526 14194 20578
rect 14590 20526 14642 20578
rect 15038 20526 15090 20578
rect 15822 20526 15874 20578
rect 16270 20526 16322 20578
rect 16606 20526 16658 20578
rect 17390 20526 17442 20578
rect 17950 20526 18002 20578
rect 18286 20526 18338 20578
rect 18734 20526 18786 20578
rect 19182 20526 19234 20578
rect 20078 20526 20130 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 1934 20190 1986 20242
rect 2718 20190 2770 20242
rect 4734 20190 4786 20242
rect 11342 20190 11394 20242
rect 18286 20190 18338 20242
rect 20526 20190 20578 20242
rect 3166 20078 3218 20130
rect 6750 20078 6802 20130
rect 10894 20078 10946 20130
rect 12462 20078 12514 20130
rect 13358 20078 13410 20130
rect 15038 20078 15090 20130
rect 20974 20078 21026 20130
rect 8542 19966 8594 20018
rect 10446 19966 10498 20018
rect 2270 19854 2322 19906
rect 4062 19854 4114 19906
rect 5182 19854 5234 19906
rect 5966 19854 6018 19906
rect 7198 19854 7250 19906
rect 7646 19854 7698 19906
rect 8206 19854 8258 19906
rect 8990 19854 9042 19906
rect 9662 19854 9714 19906
rect 12014 19854 12066 19906
rect 13022 19854 13074 19906
rect 14030 19854 14082 19906
rect 14478 19854 14530 19906
rect 15598 19854 15650 19906
rect 16046 19854 16098 19906
rect 16718 19854 16770 19906
rect 17950 19854 18002 19906
rect 18734 19854 18786 19906
rect 19294 19854 19346 19906
rect 19630 19854 19682 19906
rect 20078 19854 20130 19906
rect 21422 19854 21474 19906
rect 1710 19742 1762 19794
rect 2270 19742 2322 19794
rect 7646 19742 7698 19794
rect 8318 19742 8370 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 1822 19406 1874 19458
rect 2830 19406 2882 19458
rect 3166 19406 3218 19458
rect 5742 19406 5794 19458
rect 6190 19406 6242 19458
rect 7310 19406 7362 19458
rect 7646 19406 7698 19458
rect 9886 19406 9938 19458
rect 11342 19406 11394 19458
rect 11566 19406 11618 19458
rect 12238 19406 12290 19458
rect 12798 19406 12850 19458
rect 1934 19294 1986 19346
rect 3166 19294 3218 19346
rect 4062 19294 4114 19346
rect 5742 19294 5794 19346
rect 7086 19294 7138 19346
rect 13582 19294 13634 19346
rect 18062 19294 18114 19346
rect 19406 19294 19458 19346
rect 20302 19294 20354 19346
rect 22430 19294 22482 19346
rect 9774 19182 9826 19234
rect 10446 19182 10498 19234
rect 11678 19182 11730 19234
rect 2270 19070 2322 19122
rect 7646 19070 7698 19122
rect 8094 19070 8146 19122
rect 8990 19070 9042 19122
rect 9886 19070 9938 19122
rect 18510 19070 18562 19122
rect 18958 19070 19010 19122
rect 2718 18958 2770 19010
rect 3614 18958 3666 19010
rect 4622 18958 4674 19010
rect 5070 18958 5122 19010
rect 6302 18958 6354 19010
rect 6638 18958 6690 19010
rect 8206 18958 8258 19010
rect 8878 18958 8930 19010
rect 11230 18958 11282 19010
rect 12238 18958 12290 19010
rect 12686 18958 12738 19010
rect 14142 18958 14194 19010
rect 14702 18958 14754 19010
rect 15150 18958 15202 19010
rect 15598 18958 15650 19010
rect 15934 18958 15986 19010
rect 16606 18958 16658 19010
rect 16942 18958 16994 19010
rect 17390 18958 17442 19010
rect 19854 18958 19906 19010
rect 20750 18958 20802 19010
rect 21534 18958 21586 19010
rect 21982 18958 22034 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 3502 18622 3554 18674
rect 4846 18622 4898 18674
rect 7310 18622 7362 18674
rect 6302 18510 6354 18562
rect 6414 18510 6466 18562
rect 7198 18510 7250 18562
rect 8094 18566 8146 18618
rect 8878 18622 8930 18674
rect 9886 18622 9938 18674
rect 10894 18622 10946 18674
rect 11790 18622 11842 18674
rect 12126 18622 12178 18674
rect 12798 18622 12850 18674
rect 22430 18622 22482 18674
rect 9774 18510 9826 18562
rect 11006 18510 11058 18562
rect 12686 18510 12738 18562
rect 1822 18398 1874 18450
rect 6638 18398 6690 18450
rect 7534 18398 7586 18450
rect 7982 18398 8034 18450
rect 8654 18398 8706 18450
rect 8990 18398 9042 18450
rect 14702 18398 14754 18450
rect 17614 18398 17666 18450
rect 18174 18398 18226 18450
rect 19630 18398 19682 18450
rect 22878 18398 22930 18450
rect 2158 18286 2210 18338
rect 2718 18286 2770 18338
rect 3166 18286 3218 18338
rect 3950 18286 4002 18338
rect 4398 18286 4450 18338
rect 5294 18286 5346 18338
rect 5854 18286 5906 18338
rect 13582 18286 13634 18338
rect 14142 18286 14194 18338
rect 15150 18286 15202 18338
rect 15598 18286 15650 18338
rect 16158 18286 16210 18338
rect 16606 18286 16658 18338
rect 18622 18286 18674 18338
rect 19182 18286 19234 18338
rect 20190 18286 20242 18338
rect 20638 18286 20690 18338
rect 21086 18286 21138 18338
rect 21646 18286 21698 18338
rect 21982 18286 22034 18338
rect 3614 18174 3666 18226
rect 4398 18174 4450 18226
rect 6078 18174 6130 18226
rect 8094 18174 8146 18226
rect 9886 18174 9938 18226
rect 10894 18174 10946 18226
rect 12798 18174 12850 18226
rect 13470 18174 13522 18226
rect 14254 18174 14306 18226
rect 14590 18174 14642 18226
rect 15038 18174 15090 18226
rect 15486 18174 15538 18226
rect 16606 18174 16658 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 4062 17838 4114 17890
rect 4846 17838 4898 17890
rect 6302 17838 6354 17890
rect 8430 17838 8482 17890
rect 18958 17838 19010 17890
rect 19630 17838 19682 17890
rect 2046 17726 2098 17778
rect 3390 17726 3442 17778
rect 9102 17726 9154 17778
rect 16830 17726 16882 17778
rect 17390 17726 17442 17778
rect 18062 17726 18114 17778
rect 18958 17726 19010 17778
rect 22542 17726 22594 17778
rect 23550 17726 23602 17778
rect 2606 17614 2658 17666
rect 5630 17614 5682 17666
rect 6190 17614 6242 17666
rect 7198 17614 7250 17666
rect 7534 17614 7586 17666
rect 12014 17614 12066 17666
rect 12686 17614 12738 17666
rect 14702 17614 14754 17666
rect 15374 17614 15426 17666
rect 3950 17502 4002 17554
rect 4958 17502 5010 17554
rect 6302 17502 6354 17554
rect 8542 17502 8594 17554
rect 11230 17502 11282 17554
rect 14030 17502 14082 17554
rect 14142 17502 14194 17554
rect 3054 17390 3106 17442
rect 4846 17390 4898 17442
rect 7422 17390 7474 17442
rect 8430 17390 8482 17442
rect 12686 17390 12738 17442
rect 13806 17390 13858 17442
rect 14814 17390 14866 17442
rect 15038 17390 15090 17442
rect 16046 17390 16098 17442
rect 18510 17390 18562 17442
rect 19406 17390 19458 17442
rect 19966 17390 20018 17442
rect 20414 17390 20466 17442
rect 20862 17390 20914 17442
rect 21534 17390 21586 17442
rect 22094 17390 22146 17442
rect 23102 17390 23154 17442
rect 24334 17390 24386 17442
rect 26910 17390 26962 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 2046 17054 2098 17106
rect 2830 17054 2882 17106
rect 3054 17054 3106 17106
rect 4510 17054 4562 17106
rect 5294 17054 5346 17106
rect 6190 17054 6242 17106
rect 6974 17054 7026 17106
rect 8430 17054 8482 17106
rect 9102 17054 9154 17106
rect 9662 17054 9714 17106
rect 10334 17054 10386 17106
rect 11566 17054 11618 17106
rect 11678 17054 11730 17106
rect 13582 17054 13634 17106
rect 16494 17054 16546 17106
rect 18734 17054 18786 17106
rect 19854 17054 19906 17106
rect 22654 17054 22706 17106
rect 23550 17054 23602 17106
rect 24334 17054 24386 17106
rect 1934 16942 1986 16994
rect 2718 16942 2770 16994
rect 3726 16942 3778 16994
rect 4398 16942 4450 16994
rect 5070 16942 5122 16994
rect 5406 16942 5458 16994
rect 6414 16942 6466 16994
rect 6526 16942 6578 16994
rect 7646 16942 7698 16994
rect 8542 16942 8594 16994
rect 10222 16942 10274 16994
rect 11342 16942 11394 16994
rect 11902 16942 11954 16994
rect 12574 16942 12626 16994
rect 12686 16942 12738 16994
rect 13806 16942 13858 16994
rect 17726 16942 17778 16994
rect 18398 16942 18450 16994
rect 18510 16942 18562 16994
rect 19070 16942 19122 16994
rect 24782 16942 24834 16994
rect 27806 16942 27858 16994
rect 2270 16830 2322 16882
rect 3838 16830 3890 16882
rect 4734 16830 4786 16882
rect 7758 16830 7810 16882
rect 8206 16830 8258 16882
rect 10558 16830 10610 16882
rect 11790 16830 11842 16882
rect 14254 16830 14306 16882
rect 14590 16830 14642 16882
rect 14814 16830 14866 16882
rect 14926 16830 14978 16882
rect 15262 16830 15314 16882
rect 15710 16830 15762 16882
rect 15822 16830 15874 16882
rect 16270 16830 16322 16882
rect 16606 16830 16658 16882
rect 19742 16830 19794 16882
rect 20078 16830 20130 16882
rect 21758 16830 21810 16882
rect 26462 16830 26514 16882
rect 13694 16718 13746 16770
rect 15374 16718 15426 16770
rect 20862 16718 20914 16770
rect 21422 16718 21474 16770
rect 22206 16718 22258 16770
rect 23102 16718 23154 16770
rect 25678 16718 25730 16770
rect 26126 16718 26178 16770
rect 27022 16718 27074 16770
rect 27470 16718 27522 16770
rect 7646 16606 7698 16658
rect 12686 16606 12738 16658
rect 17838 16606 17890 16658
rect 20750 16606 20802 16658
rect 21534 16606 21586 16658
rect 27022 16606 27074 16658
rect 27694 16606 27746 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 2382 16270 2434 16322
rect 5742 16270 5794 16322
rect 6078 16270 6130 16322
rect 12798 16270 12850 16322
rect 18846 16270 18898 16322
rect 20750 16270 20802 16322
rect 4734 16158 4786 16210
rect 10558 16158 10610 16210
rect 13918 16158 13970 16210
rect 22766 16158 22818 16210
rect 23214 16158 23266 16210
rect 29486 16158 29538 16210
rect 29934 16158 29986 16210
rect 1822 16046 1874 16098
rect 2270 16046 2322 16098
rect 3054 16046 3106 16098
rect 3838 16046 3890 16098
rect 6526 16046 6578 16098
rect 7758 16046 7810 16098
rect 13694 16046 13746 16098
rect 17950 16046 18002 16098
rect 20414 16046 20466 16098
rect 21534 16046 21586 16098
rect 21870 16046 21922 16098
rect 2382 15822 2434 15874
rect 3166 15822 3218 15874
rect 3390 15822 3442 15874
rect 3950 15878 4002 15930
rect 4622 15934 4674 15986
rect 4846 15934 4898 15986
rect 5966 15934 6018 15986
rect 8430 15934 8482 15986
rect 11118 15934 11170 15986
rect 11230 15934 11282 15986
rect 11454 15934 11506 15986
rect 11902 15934 11954 15986
rect 12686 15934 12738 15986
rect 12798 15934 12850 15986
rect 14590 15934 14642 15986
rect 14702 15934 14754 15986
rect 15374 15934 15426 15986
rect 15710 15934 15762 15986
rect 16494 15934 16546 15986
rect 17166 15934 17218 15986
rect 17390 15934 17442 15986
rect 18062 15934 18114 15986
rect 18734 15934 18786 15986
rect 19406 15934 19458 15986
rect 20190 15934 20242 15986
rect 20638 15934 20690 15986
rect 4174 15822 4226 15874
rect 6862 15822 6914 15874
rect 7086 15822 7138 15874
rect 7198 15822 7250 15874
rect 12014 15822 12066 15874
rect 12238 15822 12290 15874
rect 13918 15822 13970 15874
rect 14926 15822 14978 15874
rect 16158 15822 16210 15874
rect 16382 15822 16434 15874
rect 17278 15822 17330 15874
rect 18286 15822 18338 15874
rect 19518 15822 19570 15874
rect 19742 15822 19794 15874
rect 22094 15822 22146 15874
rect 22206 15822 22258 15874
rect 22654 15822 22706 15874
rect 23998 15822 24050 15874
rect 24894 15822 24946 15874
rect 25230 15822 25282 15874
rect 26014 15822 26066 15874
rect 26462 15822 26514 15874
rect 26798 15822 26850 15874
rect 27246 15822 27298 15874
rect 27694 15822 27746 15874
rect 28254 15822 28306 15874
rect 28814 15822 28866 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 2046 15486 2098 15538
rect 2270 15486 2322 15538
rect 2830 15486 2882 15538
rect 3054 15486 3106 15538
rect 4398 15486 4450 15538
rect 5182 15486 5234 15538
rect 5406 15486 5458 15538
rect 7310 15486 7362 15538
rect 7534 15486 7586 15538
rect 8318 15486 8370 15538
rect 8430 15486 8482 15538
rect 10334 15486 10386 15538
rect 11902 15486 11954 15538
rect 12574 15486 12626 15538
rect 12798 15486 12850 15538
rect 13582 15486 13634 15538
rect 14142 15486 14194 15538
rect 16942 15486 16994 15538
rect 17838 15486 17890 15538
rect 20750 15486 20802 15538
rect 20862 15486 20914 15538
rect 21310 15486 21362 15538
rect 21534 15486 21586 15538
rect 26238 15486 26290 15538
rect 27134 15486 27186 15538
rect 30718 15486 30770 15538
rect 1934 15374 1986 15426
rect 2718 15374 2770 15426
rect 3502 15374 3554 15426
rect 3614 15374 3666 15426
rect 4286 15374 4338 15426
rect 5070 15374 5122 15426
rect 5854 15374 5906 15426
rect 6302 15374 6354 15426
rect 7086 15374 7138 15426
rect 8094 15374 8146 15426
rect 9998 15374 10050 15426
rect 10110 15374 10162 15426
rect 10894 15374 10946 15426
rect 11678 15374 11730 15426
rect 13358 15374 13410 15426
rect 18622 15374 18674 15426
rect 19742 15374 19794 15426
rect 22766 15374 22818 15426
rect 24446 15374 24498 15426
rect 24558 15374 24610 15426
rect 25678 15374 25730 15426
rect 31166 15374 31218 15426
rect 3838 15262 3890 15314
rect 4622 15262 4674 15314
rect 6078 15262 6130 15314
rect 6414 15262 6466 15314
rect 8542 15262 8594 15314
rect 8766 15262 8818 15314
rect 10782 15262 10834 15314
rect 11118 15262 11170 15314
rect 11566 15262 11618 15314
rect 12238 15262 12290 15314
rect 14590 15262 14642 15314
rect 14926 15262 14978 15314
rect 15262 15262 15314 15314
rect 15710 15262 15762 15314
rect 16158 15262 16210 15314
rect 16270 15262 16322 15314
rect 17614 15262 17666 15314
rect 17950 15262 18002 15314
rect 18510 15262 18562 15314
rect 18734 15262 18786 15314
rect 19182 15262 19234 15314
rect 19630 15262 19682 15314
rect 20302 15262 20354 15314
rect 20526 15262 20578 15314
rect 21870 15262 21922 15314
rect 22542 15262 22594 15314
rect 23214 15262 23266 15314
rect 28030 15262 28082 15314
rect 29822 15262 29874 15314
rect 7534 15150 7586 15202
rect 12462 15150 12514 15202
rect 13694 15150 13746 15202
rect 14814 15150 14866 15202
rect 15934 15150 15986 15202
rect 22990 15150 23042 15202
rect 23774 15150 23826 15202
rect 25790 15150 25842 15202
rect 26798 15150 26850 15202
rect 27582 15150 27634 15202
rect 28590 15150 28642 15202
rect 29038 15150 29090 15202
rect 29486 15150 29538 15202
rect 30382 15150 30434 15202
rect 31726 15150 31778 15202
rect 32174 15150 32226 15202
rect 32622 15150 32674 15202
rect 21198 15038 21250 15090
rect 23662 15038 23714 15090
rect 24446 15038 24498 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16270 14702 16322 14754
rect 17390 14702 17442 14754
rect 19406 14702 19458 14754
rect 31950 14702 32002 14754
rect 33518 14702 33570 14754
rect 2158 14590 2210 14642
rect 8766 14590 8818 14642
rect 12238 14590 12290 14642
rect 14814 14590 14866 14642
rect 23774 14590 23826 14642
rect 25902 14590 25954 14642
rect 27470 14590 27522 14642
rect 28030 14590 28082 14642
rect 2382 14478 2434 14530
rect 3838 14478 3890 14530
rect 6078 14478 6130 14530
rect 8206 14478 8258 14530
rect 11566 14478 11618 14530
rect 12686 14478 12738 14530
rect 13022 14478 13074 14530
rect 14030 14478 14082 14530
rect 15038 14478 15090 14530
rect 16270 14478 16322 14530
rect 16830 14478 16882 14530
rect 17054 14478 17106 14530
rect 18398 14478 18450 14530
rect 19518 14478 19570 14530
rect 20078 14478 20130 14530
rect 21646 14478 21698 14530
rect 22990 14478 23042 14530
rect 27022 14478 27074 14530
rect 3502 14366 3554 14418
rect 4286 14366 4338 14418
rect 7198 14366 7250 14418
rect 10894 14366 10946 14418
rect 12798 14366 12850 14418
rect 14142 14366 14194 14418
rect 15934 14366 15986 14418
rect 18062 14366 18114 14418
rect 20526 14366 20578 14418
rect 21982 14366 22034 14418
rect 33294 14366 33346 14418
rect 2942 14254 2994 14306
rect 3614 14254 3666 14306
rect 4398 14254 4450 14306
rect 5854 14254 5906 14306
rect 5966 14254 6018 14306
rect 6750 14254 6802 14306
rect 7310 14254 7362 14306
rect 7534 14254 7586 14306
rect 7870 14254 7922 14306
rect 8094 14254 8146 14306
rect 14366 14254 14418 14306
rect 15374 14254 15426 14306
rect 17278 14254 17330 14306
rect 18174 14254 18226 14306
rect 19406 14254 19458 14306
rect 20302 14254 20354 14306
rect 20638 14254 20690 14306
rect 22094 14254 22146 14306
rect 22206 14254 22258 14306
rect 26350 14254 26402 14306
rect 26462 14254 26514 14306
rect 26686 14254 26738 14306
rect 27582 14254 27634 14306
rect 28478 14254 28530 14306
rect 29598 14254 29650 14306
rect 29934 14254 29986 14306
rect 30382 14254 30434 14306
rect 30942 14254 30994 14306
rect 31614 14254 31666 14306
rect 32062 14254 32114 14306
rect 32398 14254 32450 14306
rect 32846 14254 32898 14306
rect 33854 14254 33906 14306
rect 34302 14254 34354 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 8094 13918 8146 13970
rect 8878 13918 8930 13970
rect 10110 13918 10162 13970
rect 10222 13918 10274 13970
rect 10334 13918 10386 13970
rect 11118 13918 11170 13970
rect 11790 13918 11842 13970
rect 12014 13918 12066 13970
rect 12574 13918 12626 13970
rect 13582 13918 13634 13970
rect 14590 13918 14642 13970
rect 17054 13918 17106 13970
rect 19070 13918 19122 13970
rect 6414 13806 6466 13858
rect 7086 13806 7138 13858
rect 7310 13806 7362 13858
rect 8206 13806 8258 13858
rect 8766 13806 8818 13858
rect 12462 13806 12514 13858
rect 12798 13806 12850 13858
rect 13246 13806 13298 13858
rect 13358 13806 13410 13858
rect 14366 13806 14418 13858
rect 14814 13806 14866 13858
rect 15374 13806 15426 13858
rect 15822 13806 15874 13858
rect 16830 13806 16882 13858
rect 18062 13806 18114 13858
rect 18734 13806 18786 13858
rect 18846 13806 18898 13858
rect 19518 13806 19570 13858
rect 19630 13862 19682 13914
rect 20190 13918 20242 13970
rect 20414 13918 20466 13970
rect 21646 13918 21698 13970
rect 21758 13918 21810 13970
rect 24558 13918 24610 13970
rect 28142 13918 28194 13970
rect 32174 13918 32226 13970
rect 23326 13806 23378 13858
rect 24446 13806 24498 13858
rect 27358 13806 27410 13858
rect 4846 13694 4898 13746
rect 5518 13694 5570 13746
rect 6302 13694 6354 13746
rect 7870 13694 7922 13746
rect 9102 13694 9154 13746
rect 9886 13694 9938 13746
rect 10446 13694 10498 13746
rect 11678 13694 11730 13746
rect 15598 13694 15650 13746
rect 16718 13694 16770 13746
rect 17950 13694 18002 13746
rect 19854 13694 19906 13746
rect 20526 13694 20578 13746
rect 21534 13694 21586 13746
rect 22206 13694 22258 13746
rect 23550 13694 23602 13746
rect 26014 13694 26066 13746
rect 26350 13694 26402 13746
rect 26686 13694 26738 13746
rect 27134 13694 27186 13746
rect 27470 13694 27522 13746
rect 27918 13694 27970 13746
rect 28254 13694 28306 13746
rect 29822 13694 29874 13746
rect 1934 13582 1986 13634
rect 4062 13582 4114 13634
rect 5742 13582 5794 13634
rect 7422 13582 7474 13634
rect 15486 13582 15538 13634
rect 20974 13582 21026 13634
rect 22654 13582 22706 13634
rect 22766 13582 22818 13634
rect 25566 13582 25618 13634
rect 26238 13582 26290 13634
rect 28814 13582 28866 13634
rect 29374 13582 29426 13634
rect 30270 13582 30322 13634
rect 30718 13582 30770 13634
rect 31166 13582 31218 13634
rect 31726 13582 31778 13634
rect 32622 13582 32674 13634
rect 33518 13582 33570 13634
rect 34078 13582 34130 13634
rect 34526 13582 34578 13634
rect 34862 13582 34914 13634
rect 35422 13582 35474 13634
rect 35870 13582 35922 13634
rect 6414 13470 6466 13522
rect 14478 13470 14530 13522
rect 18062 13470 18114 13522
rect 23886 13470 23938 13522
rect 24558 13470 24610 13522
rect 28926 13470 28978 13522
rect 29598 13470 29650 13522
rect 30270 13470 30322 13522
rect 33630 13470 33682 13522
rect 34862 13470 34914 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 4622 13134 4674 13186
rect 6078 13134 6130 13186
rect 14366 13134 14418 13186
rect 14926 13134 14978 13186
rect 25566 13134 25618 13186
rect 27470 13134 27522 13186
rect 33518 13134 33570 13186
rect 35982 13134 36034 13186
rect 3950 13022 4002 13074
rect 7310 13022 7362 13074
rect 8206 13022 8258 13074
rect 9662 13022 9714 13074
rect 24446 13022 24498 13074
rect 33742 13022 33794 13074
rect 2046 12910 2098 12962
rect 3166 12910 3218 12962
rect 5742 12910 5794 12962
rect 5966 12910 6018 12962
rect 8430 12910 8482 12962
rect 12574 12910 12626 12962
rect 14590 12910 14642 12962
rect 14814 12910 14866 12962
rect 15710 12910 15762 12962
rect 15822 12910 15874 12962
rect 16270 12910 16322 12962
rect 16606 12910 16658 12962
rect 18958 12910 19010 12962
rect 19294 12910 19346 12962
rect 20078 12910 20130 12962
rect 20414 12910 20466 12962
rect 23326 12910 23378 12962
rect 23550 12910 23602 12962
rect 24670 12910 24722 12962
rect 26238 12910 26290 12962
rect 26462 12910 26514 12962
rect 26910 12910 26962 12962
rect 32846 12910 32898 12962
rect 2270 12798 2322 12850
rect 4062 12798 4114 12850
rect 6974 12798 7026 12850
rect 11790 12798 11842 12850
rect 13694 12798 13746 12850
rect 14254 12798 14306 12850
rect 17166 12798 17218 12850
rect 17390 12798 17442 12850
rect 17614 12798 17666 12850
rect 17726 12798 17778 12850
rect 19742 12798 19794 12850
rect 21870 12798 21922 12850
rect 22542 12798 22594 12850
rect 22654 12798 22706 12850
rect 23774 12798 23826 12850
rect 25678 12798 25730 12850
rect 27358 12798 27410 12850
rect 27470 12798 27522 12850
rect 28254 12798 28306 12850
rect 28366 12798 28418 12850
rect 29598 12798 29650 12850
rect 30270 12798 30322 12850
rect 30942 12798 30994 12850
rect 31726 12798 31778 12850
rect 32286 12798 32338 12850
rect 35534 12798 35586 12850
rect 3054 12686 3106 12738
rect 3838 12686 3890 12738
rect 4734 12686 4786 12738
rect 4846 12686 4898 12738
rect 7198 12686 7250 12738
rect 7422 12686 7474 12738
rect 7534 12686 7586 12738
rect 8766 12686 8818 12738
rect 15934 12686 15986 12738
rect 16942 12686 16994 12738
rect 17278 12686 17330 12738
rect 17838 12686 17890 12738
rect 19070 12686 19122 12738
rect 20190 12686 20242 12738
rect 20862 12686 20914 12738
rect 21534 12686 21586 12738
rect 21758 12686 21810 12738
rect 22318 12686 22370 12738
rect 23886 12686 23938 12738
rect 25006 12686 25058 12738
rect 26350 12686 26402 12738
rect 28030 12686 28082 12738
rect 28814 12686 28866 12738
rect 29710 12686 29762 12738
rect 30382 12686 30434 12738
rect 31054 12686 31106 12738
rect 31614 12686 31666 12738
rect 32398 12686 32450 12738
rect 33294 12686 33346 12738
rect 34190 12686 34242 12738
rect 34750 12686 34802 12738
rect 35086 12686 35138 12738
rect 35982 12686 36034 12738
rect 36430 12686 36482 12738
rect 37438 12686 37490 12738
rect 37886 12686 37938 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 1934 12350 1986 12402
rect 2606 12350 2658 12402
rect 3726 12350 3778 12402
rect 4622 12350 4674 12402
rect 5406 12350 5458 12402
rect 6750 12350 6802 12402
rect 6974 12350 7026 12402
rect 8206 12350 8258 12402
rect 8430 12350 8482 12402
rect 9102 12350 9154 12402
rect 17614 12350 17666 12402
rect 18846 12350 18898 12402
rect 23214 12350 23266 12402
rect 24222 12350 24274 12402
rect 25566 12350 25618 12402
rect 25790 12350 25842 12402
rect 33518 12350 33570 12402
rect 34862 12350 34914 12402
rect 36542 12350 36594 12402
rect 40462 12350 40514 12402
rect 41470 12350 41522 12402
rect 42030 12350 42082 12402
rect 1822 12238 1874 12290
rect 2494 12238 2546 12290
rect 3950 12238 4002 12290
rect 4510 12238 4562 12290
rect 5182 12238 5234 12290
rect 5630 12238 5682 12290
rect 11006 12238 11058 12290
rect 17838 12238 17890 12290
rect 17950 12238 18002 12290
rect 18622 12238 18674 12290
rect 20302 12238 20354 12290
rect 23102 12238 23154 12290
rect 23662 12238 23714 12290
rect 25902 12238 25954 12290
rect 27470 12238 27522 12290
rect 30270 12238 30322 12290
rect 32734 12238 32786 12290
rect 33966 12238 34018 12290
rect 2830 12126 2882 12178
rect 3502 12126 3554 12178
rect 3726 12126 3778 12178
rect 7422 12126 7474 12178
rect 7982 12126 8034 12178
rect 9774 12126 9826 12178
rect 16718 12126 16770 12178
rect 18510 12126 18562 12178
rect 19630 12126 19682 12178
rect 23326 12126 23378 12178
rect 23438 12126 23490 12178
rect 24558 12126 24610 12178
rect 26686 12126 26738 12178
rect 30158 12126 30210 12178
rect 32846 12126 32898 12178
rect 6302 12014 6354 12066
rect 6862 12014 6914 12066
rect 8094 12014 8146 12066
rect 10222 12014 10274 12066
rect 14590 12014 14642 12066
rect 22430 12014 22482 12066
rect 24782 12014 24834 12066
rect 29598 12014 29650 12066
rect 30942 12014 30994 12066
rect 31614 12014 31666 12066
rect 32062 12014 32114 12066
rect 34414 12014 34466 12066
rect 35646 12014 35698 12066
rect 36094 12014 36146 12066
rect 36990 12014 37042 12066
rect 37886 12014 37938 12066
rect 37998 12014 38050 12066
rect 38558 12014 38610 12066
rect 38894 12014 38946 12066
rect 39566 12014 39618 12066
rect 5742 11902 5794 11954
rect 10894 11902 10946 11954
rect 30830 11902 30882 11954
rect 31502 11902 31554 11954
rect 32734 11902 32786 11954
rect 33518 11902 33570 11954
rect 33854 11902 33906 11954
rect 34414 11902 34466 11954
rect 35534 11902 35586 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 9326 11566 9378 11618
rect 10782 11566 10834 11618
rect 15934 11566 15986 11618
rect 40798 11566 40850 11618
rect 41694 11566 41746 11618
rect 1822 11454 1874 11506
rect 7310 11454 7362 11506
rect 8990 11454 9042 11506
rect 12574 11454 12626 11506
rect 14030 11454 14082 11506
rect 18174 11454 18226 11506
rect 21870 11454 21922 11506
rect 27918 11454 27970 11506
rect 36766 11454 36818 11506
rect 41694 11454 41746 11506
rect 4734 11342 4786 11394
rect 5742 11342 5794 11394
rect 6078 11342 6130 11394
rect 6190 11342 6242 11394
rect 6414 11342 6466 11394
rect 6638 11342 6690 11394
rect 7086 11342 7138 11394
rect 7534 11342 7586 11394
rect 8878 11342 8930 11394
rect 9102 11342 9154 11394
rect 9550 11342 9602 11394
rect 9774 11342 9826 11394
rect 10222 11342 10274 11394
rect 10558 11342 10610 11394
rect 11006 11342 11058 11394
rect 11230 11342 11282 11394
rect 12238 11342 12290 11394
rect 12686 11342 12738 11394
rect 12910 11342 12962 11394
rect 17390 11342 17442 11394
rect 19406 11342 19458 11394
rect 20414 11342 20466 11394
rect 21646 11342 21698 11394
rect 22206 11342 22258 11394
rect 23550 11342 23602 11394
rect 23886 11342 23938 11394
rect 23998 11342 24050 11394
rect 24558 11342 24610 11394
rect 25678 11342 25730 11394
rect 26014 11342 26066 11394
rect 26686 11342 26738 11394
rect 28366 11342 28418 11394
rect 28702 11342 28754 11394
rect 29934 11342 29986 11394
rect 30606 11342 30658 11394
rect 31726 11342 31778 11394
rect 33182 11342 33234 11394
rect 33854 11342 33906 11394
rect 37662 11342 37714 11394
rect 37886 11342 37938 11394
rect 37998 11342 38050 11394
rect 38670 11342 38722 11394
rect 39006 11342 39058 11394
rect 39230 11342 39282 11394
rect 3950 11230 4002 11282
rect 7758 11230 7810 11282
rect 13694 11230 13746 11282
rect 14702 11230 14754 11282
rect 16158 11230 16210 11282
rect 17502 11230 17554 11282
rect 18622 11230 18674 11282
rect 24894 11230 24946 11282
rect 25790 11230 25842 11282
rect 27470 11230 27522 11282
rect 29598 11230 29650 11282
rect 31054 11230 31106 11282
rect 31838 11230 31890 11282
rect 32510 11230 32562 11282
rect 32622 11230 32674 11282
rect 34638 11230 34690 11282
rect 37550 11230 37602 11282
rect 6078 11118 6130 11170
rect 8318 11118 8370 11170
rect 10670 11118 10722 11170
rect 11678 11118 11730 11170
rect 12462 11118 12514 11170
rect 14814 11118 14866 11170
rect 15598 11118 15650 11170
rect 17166 11118 17218 11170
rect 17614 11118 17666 11170
rect 18734 11118 18786 11170
rect 18958 11118 19010 11170
rect 19630 11118 19682 11170
rect 19854 11118 19906 11170
rect 19966 11118 20018 11170
rect 20638 11118 20690 11170
rect 20862 11118 20914 11170
rect 20974 11118 21026 11170
rect 21870 11118 21922 11170
rect 22094 11118 22146 11170
rect 22766 11118 22818 11170
rect 23662 11118 23714 11170
rect 23774 11118 23826 11170
rect 24782 11118 24834 11170
rect 26350 11118 26402 11170
rect 26574 11118 26626 11170
rect 27134 11118 27186 11170
rect 27358 11118 27410 11170
rect 28590 11118 28642 11170
rect 29710 11118 29762 11170
rect 30270 11118 30322 11170
rect 30494 11118 30546 11170
rect 32062 11118 32114 11170
rect 32846 11118 32898 11170
rect 39678 11118 39730 11170
rect 40350 11118 40402 11170
rect 40798 11118 40850 11170
rect 41246 11118 41298 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4174 10782 4226 10834
rect 4286 10782 4338 10834
rect 4398 10782 4450 10834
rect 4510 10782 4562 10834
rect 6638 10782 6690 10834
rect 7422 10782 7474 10834
rect 8430 10782 8482 10834
rect 9662 10782 9714 10834
rect 15486 10782 15538 10834
rect 15710 10782 15762 10834
rect 16270 10782 16322 10834
rect 16382 10782 16434 10834
rect 17614 10782 17666 10834
rect 32846 10782 32898 10834
rect 34862 10782 34914 10834
rect 35422 10782 35474 10834
rect 36094 10782 36146 10834
rect 38222 10782 38274 10834
rect 40574 10782 40626 10834
rect 41470 10782 41522 10834
rect 1934 10670 1986 10722
rect 5182 10670 5234 10722
rect 5630 10670 5682 10722
rect 7198 10670 7250 10722
rect 7534 10670 7586 10722
rect 10670 10670 10722 10722
rect 15374 10670 15426 10722
rect 16494 10670 16546 10722
rect 17054 10670 17106 10722
rect 17838 10670 17890 10722
rect 33966 10670 34018 10722
rect 36206 10670 36258 10722
rect 36878 10670 36930 10722
rect 3950 10558 4002 10610
rect 5406 10558 5458 10610
rect 6190 10558 6242 10610
rect 6414 10558 6466 10610
rect 7758 10558 7810 10610
rect 9774 10558 9826 10610
rect 9998 10558 10050 10610
rect 10334 10558 10386 10610
rect 11230 10558 11282 10610
rect 14702 10558 14754 10610
rect 17950 10558 18002 10610
rect 18510 10558 18562 10610
rect 24222 10558 24274 10610
rect 24558 10558 24610 10610
rect 24894 10558 24946 10610
rect 26014 10558 26066 10610
rect 29598 10558 29650 10610
rect 33518 10558 33570 10610
rect 34190 10558 34242 10610
rect 34750 10558 34802 10610
rect 35870 10558 35922 10610
rect 36990 10558 37042 10610
rect 37998 10558 38050 10610
rect 40126 10558 40178 10610
rect 3278 10446 3330 10498
rect 6750 10446 6802 10498
rect 8990 10446 9042 10498
rect 11902 10446 11954 10498
rect 14030 10446 14082 10498
rect 20526 10446 20578 10498
rect 24446 10446 24498 10498
rect 26798 10446 26850 10498
rect 28926 10446 28978 10498
rect 30270 10446 30322 10498
rect 32398 10446 32450 10498
rect 33742 10446 33794 10498
rect 37438 10446 37490 10498
rect 38222 10446 38274 10498
rect 38782 10446 38834 10498
rect 39230 10446 39282 10498
rect 39678 10446 39730 10498
rect 41918 10446 41970 10498
rect 5294 10334 5346 10386
rect 10222 10334 10274 10386
rect 11342 10334 11394 10386
rect 34862 10334 34914 10386
rect 36878 10334 36930 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 4958 9998 5010 10050
rect 7310 9998 7362 10050
rect 10110 9998 10162 10050
rect 17166 9998 17218 10050
rect 27358 9998 27410 10050
rect 27806 9998 27858 10050
rect 2158 9886 2210 9938
rect 2718 9886 2770 9938
rect 3054 9886 3106 9938
rect 4846 9886 4898 9938
rect 6414 9886 6466 9938
rect 14030 9886 14082 9938
rect 16046 9886 16098 9938
rect 18510 9886 18562 9938
rect 21870 9886 21922 9938
rect 22878 9886 22930 9938
rect 24110 9886 24162 9938
rect 26238 9886 26290 9938
rect 26686 9886 26738 9938
rect 27470 9886 27522 9938
rect 27694 9886 27746 9938
rect 28478 9886 28530 9938
rect 30158 9886 30210 9938
rect 33294 9886 33346 9938
rect 35422 9886 35474 9938
rect 37662 9886 37714 9938
rect 38670 9886 38722 9938
rect 40574 9886 40626 9938
rect 41470 9886 41522 9938
rect 41918 9886 41970 9938
rect 3838 9774 3890 9826
rect 4062 9774 4114 9826
rect 6190 9774 6242 9826
rect 7646 9774 7698 9826
rect 9774 9774 9826 9826
rect 10222 9774 10274 9826
rect 11566 9774 11618 9826
rect 13694 9774 13746 9826
rect 13918 9774 13970 9826
rect 14142 9774 14194 9826
rect 14366 9774 14418 9826
rect 16158 9774 16210 9826
rect 17726 9774 17778 9826
rect 18622 9774 18674 9826
rect 18846 9774 18898 9826
rect 20638 9774 20690 9826
rect 20862 9774 20914 9826
rect 22430 9774 22482 9826
rect 23438 9774 23490 9826
rect 29822 9774 29874 9826
rect 30046 9774 30098 9826
rect 30382 9774 30434 9826
rect 31838 9774 31890 9826
rect 32510 9774 32562 9826
rect 36206 9774 36258 9826
rect 37886 9774 37938 9826
rect 38110 9774 38162 9826
rect 40126 9774 40178 9826
rect 41022 9774 41074 9826
rect 1822 9662 1874 9714
rect 2046 9662 2098 9714
rect 3614 9662 3666 9714
rect 5742 9662 5794 9714
rect 5966 9662 6018 9714
rect 6638 9662 6690 9714
rect 7870 9662 7922 9714
rect 8990 9662 9042 9714
rect 9550 9662 9602 9714
rect 10782 9662 10834 9714
rect 12126 9662 12178 9714
rect 12686 9662 12738 9714
rect 12798 9662 12850 9714
rect 14926 9662 14978 9714
rect 16830 9662 16882 9714
rect 17838 9662 17890 9714
rect 18398 9662 18450 9714
rect 19518 9662 19570 9714
rect 19630 9662 19682 9714
rect 19854 9662 19906 9714
rect 20302 9662 20354 9714
rect 28814 9662 28866 9714
rect 31166 9662 31218 9714
rect 31502 9662 31554 9714
rect 37550 9662 37602 9714
rect 38782 9662 38834 9714
rect 39006 9662 39058 9714
rect 39566 9662 39618 9714
rect 2942 9550 2994 9602
rect 3950 9550 4002 9602
rect 4174 9550 4226 9602
rect 6526 9550 6578 9602
rect 8430 9550 8482 9602
rect 9998 9550 10050 9602
rect 10894 9550 10946 9602
rect 11118 9550 11170 9602
rect 13022 9550 13074 9602
rect 15038 9550 15090 9602
rect 17054 9550 17106 9602
rect 20526 9550 20578 9602
rect 21758 9550 21810 9602
rect 21982 9550 22034 9602
rect 28590 9550 28642 9602
rect 31838 9550 31890 9602
rect 35870 9550 35922 9602
rect 36094 9550 36146 9602
rect 36654 9550 36706 9602
rect 39678 9550 39730 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 5406 9214 5458 9266
rect 6526 9214 6578 9266
rect 7086 9214 7138 9266
rect 7198 9214 7250 9266
rect 9998 9214 10050 9266
rect 10110 9214 10162 9266
rect 11678 9214 11730 9266
rect 13470 9214 13522 9266
rect 14702 9214 14754 9266
rect 15262 9214 15314 9266
rect 16158 9214 16210 9266
rect 16270 9214 16322 9266
rect 17838 9214 17890 9266
rect 19182 9214 19234 9266
rect 19294 9214 19346 9266
rect 20414 9214 20466 9266
rect 20638 9214 20690 9266
rect 32062 9214 32114 9266
rect 32622 9214 32674 9266
rect 33518 9214 33570 9266
rect 33742 9214 33794 9266
rect 39230 9214 39282 9266
rect 39790 9214 39842 9266
rect 40238 9214 40290 9266
rect 41470 9214 41522 9266
rect 41918 9214 41970 9266
rect 3950 9102 4002 9154
rect 6414 9102 6466 9154
rect 7534 9102 7586 9154
rect 8318 9102 8370 9154
rect 8766 9102 8818 9154
rect 11118 9102 11170 9154
rect 12238 9102 12290 9154
rect 13358 9102 13410 9154
rect 14030 9102 14082 9154
rect 16718 9102 16770 9154
rect 18062 9102 18114 9154
rect 18286 9102 18338 9154
rect 29486 9102 29538 9154
rect 30270 9102 30322 9154
rect 31278 9102 31330 9154
rect 35422 9102 35474 9154
rect 38110 9102 38162 9154
rect 4734 8990 4786 9042
rect 5854 8990 5906 9042
rect 6302 8990 6354 9042
rect 7310 8990 7362 9042
rect 8542 8990 8594 9042
rect 9886 8990 9938 9042
rect 10446 8990 10498 9042
rect 12686 8990 12738 9042
rect 14254 8990 14306 9042
rect 15486 8990 15538 9042
rect 15822 8990 15874 9042
rect 16494 8990 16546 9042
rect 17614 8990 17666 9042
rect 20862 8990 20914 9042
rect 21422 8990 21474 9042
rect 22094 8990 22146 9042
rect 28590 8990 28642 9042
rect 29262 8990 29314 9042
rect 30942 8990 30994 9042
rect 33854 8990 33906 9042
rect 34750 8990 34802 9042
rect 38222 8990 38274 9042
rect 38446 8990 38498 9042
rect 38670 8990 38722 9042
rect 1822 8878 1874 8930
rect 5294 8878 5346 8930
rect 13582 8878 13634 8930
rect 15374 8878 15426 8930
rect 19854 8878 19906 8930
rect 20750 8878 20802 8930
rect 22766 8878 22818 8930
rect 24894 8878 24946 8930
rect 25678 8878 25730 8930
rect 27806 8878 27858 8930
rect 30270 8878 30322 8930
rect 31838 8878 31890 8930
rect 37550 8878 37602 8930
rect 39342 8878 39394 8930
rect 40686 8878 40738 8930
rect 8206 8766 8258 8818
rect 13806 8766 13858 8818
rect 19406 8766 19458 8818
rect 30046 8766 30098 8818
rect 30942 8766 30994 8818
rect 32174 8766 32226 8818
rect 32398 8766 32450 8818
rect 33070 8766 33122 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 1934 8430 1986 8482
rect 14142 8430 14194 8482
rect 15262 8430 15314 8482
rect 35534 8430 35586 8482
rect 37550 8430 37602 8482
rect 1822 8318 1874 8370
rect 3054 8318 3106 8370
rect 5966 8318 6018 8370
rect 7086 8318 7138 8370
rect 8206 8318 8258 8370
rect 12798 8318 12850 8370
rect 13806 8318 13858 8370
rect 15150 8318 15202 8370
rect 15822 8318 15874 8370
rect 20526 8318 20578 8370
rect 21982 8318 22034 8370
rect 31054 8318 31106 8370
rect 31166 8318 31218 8370
rect 31838 8318 31890 8370
rect 34526 8318 34578 8370
rect 39566 8318 39618 8370
rect 40126 8318 40178 8370
rect 41582 8318 41634 8370
rect 2494 8206 2546 8258
rect 2718 8206 2770 8258
rect 3950 8206 4002 8258
rect 6190 8206 6242 8258
rect 6302 8206 6354 8258
rect 9326 8206 9378 8258
rect 9998 8206 10050 8258
rect 13918 8206 13970 8258
rect 14366 8206 14418 8258
rect 14702 8206 14754 8258
rect 16046 8206 16098 8258
rect 17166 8206 17218 8258
rect 17614 8206 17666 8258
rect 19294 8206 19346 8258
rect 19518 8206 19570 8258
rect 20302 8206 20354 8258
rect 22206 8206 22258 8258
rect 23102 8206 23154 8258
rect 29822 8206 29874 8258
rect 30382 8206 30434 8258
rect 31390 8206 31442 8258
rect 32510 8206 32562 8258
rect 35646 8206 35698 8258
rect 36206 8206 36258 8258
rect 36542 8206 36594 8258
rect 38670 8206 38722 8258
rect 39230 8206 39282 8258
rect 2942 8094 2994 8146
rect 3502 8094 3554 8146
rect 4734 8094 4786 8146
rect 5070 8094 5122 8146
rect 5742 8094 5794 8146
rect 6638 8094 6690 8146
rect 10670 8094 10722 8146
rect 13694 8094 13746 8146
rect 16942 8094 16994 8146
rect 18846 8094 18898 8146
rect 19070 8094 19122 8146
rect 19742 8094 19794 8146
rect 20862 8094 20914 8146
rect 21870 8094 21922 8146
rect 22430 8094 22482 8146
rect 26798 8094 26850 8146
rect 33966 8094 34018 8146
rect 34638 8094 34690 8146
rect 34750 8094 34802 8146
rect 38558 8094 38610 8146
rect 40238 8094 40290 8146
rect 41134 8094 41186 8146
rect 3726 7982 3778 8034
rect 3838 7982 3890 8034
rect 4062 7982 4114 8034
rect 4846 7982 4898 8034
rect 5630 7982 5682 8034
rect 7646 7982 7698 8034
rect 8766 7982 8818 8034
rect 8878 7982 8930 8034
rect 8990 7982 9042 8034
rect 16382 7982 16434 8034
rect 17278 7982 17330 8034
rect 17390 7982 17442 8034
rect 18286 7982 18338 8034
rect 19854 7982 19906 8034
rect 20638 7982 20690 8034
rect 28702 7982 28754 8034
rect 30270 7982 30322 8034
rect 30494 7982 30546 8034
rect 32622 7982 32674 8034
rect 32734 7982 32786 8034
rect 32958 7982 33010 8034
rect 33742 7982 33794 8034
rect 33854 7982 33906 8034
rect 35534 7982 35586 8034
rect 36318 7982 36370 8034
rect 37662 7982 37714 8034
rect 37774 7982 37826 8034
rect 38334 7982 38386 8034
rect 39454 7982 39506 8034
rect 40686 7982 40738 8034
rect 42030 7982 42082 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 7086 7646 7138 7698
rect 7310 7646 7362 7698
rect 9102 7646 9154 7698
rect 10782 7646 10834 7698
rect 11006 7646 11058 7698
rect 17614 7646 17666 7698
rect 17726 7646 17778 7698
rect 17950 7646 18002 7698
rect 20302 7646 20354 7698
rect 24446 7646 24498 7698
rect 25790 7646 25842 7698
rect 27582 7646 27634 7698
rect 27694 7646 27746 7698
rect 27806 7646 27858 7698
rect 38334 7646 38386 7698
rect 41806 7646 41858 7698
rect 3950 7534 4002 7586
rect 7982 7534 8034 7586
rect 10446 7534 10498 7586
rect 13134 7534 13186 7586
rect 18174 7534 18226 7586
rect 25902 7534 25954 7586
rect 29150 7534 29202 7586
rect 31950 7534 32002 7586
rect 32286 7534 32338 7586
rect 32510 7534 32562 7586
rect 33630 7534 33682 7586
rect 33854 7534 33906 7586
rect 35534 7534 35586 7586
rect 38222 7534 38274 7586
rect 4734 7422 4786 7474
rect 5518 7422 5570 7474
rect 6190 7422 6242 7474
rect 6862 7422 6914 7474
rect 6974 7422 7026 7474
rect 8206 7422 8258 7474
rect 8430 7422 8482 7474
rect 10558 7422 10610 7474
rect 16606 7422 16658 7474
rect 18734 7422 18786 7474
rect 19070 7422 19122 7474
rect 19630 7422 19682 7474
rect 20862 7422 20914 7474
rect 24222 7422 24274 7474
rect 27134 7422 27186 7474
rect 28478 7422 28530 7474
rect 34750 7422 34802 7474
rect 40126 7422 40178 7474
rect 1822 7310 1874 7362
rect 5966 7310 6018 7362
rect 9774 7310 9826 7362
rect 10670 7310 10722 7362
rect 19406 7310 19458 7362
rect 19518 7310 19570 7362
rect 21534 7310 21586 7362
rect 23662 7310 23714 7362
rect 26686 7310 26738 7362
rect 31278 7310 31330 7362
rect 32062 7310 32114 7362
rect 33966 7310 34018 7362
rect 37662 7310 37714 7362
rect 39230 7310 39282 7362
rect 40686 7310 40738 7362
rect 41694 7310 41746 7362
rect 5406 7198 5458 7250
rect 5742 7198 5794 7250
rect 8654 7198 8706 7250
rect 19182 7198 19234 7250
rect 24558 7198 24610 7250
rect 25678 7198 25730 7250
rect 26574 7198 26626 7250
rect 40798 7198 40850 7250
rect 41582 7198 41634 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 15598 6862 15650 6914
rect 17054 6862 17106 6914
rect 28702 6862 28754 6914
rect 28926 6862 28978 6914
rect 29598 6862 29650 6914
rect 29934 6862 29986 6914
rect 36318 6862 36370 6914
rect 4174 6750 4226 6802
rect 5966 6750 6018 6802
rect 7422 6750 7474 6802
rect 11566 6750 11618 6802
rect 15262 6750 15314 6802
rect 20526 6750 20578 6802
rect 23550 6750 23602 6802
rect 31950 6750 32002 6802
rect 34078 6750 34130 6802
rect 36094 6750 36146 6802
rect 36766 6750 36818 6802
rect 37774 6750 37826 6802
rect 41246 6750 41298 6802
rect 4734 6638 4786 6690
rect 6190 6638 6242 6690
rect 6414 6638 6466 6690
rect 6638 6638 6690 6690
rect 7534 6638 7586 6690
rect 9550 6638 9602 6690
rect 9998 6638 10050 6690
rect 10334 6638 10386 6690
rect 10446 6638 10498 6690
rect 10558 6638 10610 6690
rect 12238 6638 12290 6690
rect 12686 6638 12738 6690
rect 14366 6638 14418 6690
rect 15150 6638 15202 6690
rect 15374 6638 15426 6690
rect 15710 6638 15762 6690
rect 16494 6638 16546 6690
rect 17278 6638 17330 6690
rect 18622 6638 18674 6690
rect 18846 6638 18898 6690
rect 20190 6638 20242 6690
rect 20414 6638 20466 6690
rect 20750 6638 20802 6690
rect 22318 6638 22370 6690
rect 28254 6638 28306 6690
rect 30606 6638 30658 6690
rect 31166 6638 31218 6690
rect 34862 6638 34914 6690
rect 35086 6638 35138 6690
rect 35534 6638 35586 6690
rect 35982 6638 36034 6690
rect 37886 6638 37938 6690
rect 40126 6638 40178 6690
rect 40798 6638 40850 6690
rect 41918 6638 41970 6690
rect 2158 6526 2210 6578
rect 2830 6526 2882 6578
rect 5742 6526 5794 6578
rect 7870 6526 7922 6578
rect 8430 6526 8482 6578
rect 9214 6526 9266 6578
rect 9326 6526 9378 6578
rect 12462 6526 12514 6578
rect 13806 6526 13858 6578
rect 14142 6526 14194 6578
rect 16046 6526 16098 6578
rect 16830 6526 16882 6578
rect 17502 6526 17554 6578
rect 18398 6526 18450 6578
rect 19070 6526 19122 6578
rect 19294 6526 19346 6578
rect 30494 6526 30546 6578
rect 38110 6526 38162 6578
rect 39006 6526 39058 6578
rect 2046 6414 2098 6466
rect 4846 6414 4898 6466
rect 5070 6414 5122 6466
rect 5630 6414 5682 6466
rect 11118 6414 11170 6466
rect 12574 6414 12626 6466
rect 12798 6414 12850 6466
rect 16942 6414 16994 6466
rect 18286 6414 18338 6466
rect 20638 6414 20690 6466
rect 21646 6414 21698 6466
rect 21758 6414 21810 6466
rect 21870 6414 21922 6466
rect 28702 6414 28754 6466
rect 29822 6414 29874 6466
rect 35310 6414 35362 6466
rect 37662 6414 37714 6466
rect 42030 6414 42082 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 10334 6078 10386 6130
rect 16942 6078 16994 6130
rect 23774 6078 23826 6130
rect 24446 6078 24498 6130
rect 24782 6078 24834 6130
rect 26798 6078 26850 6130
rect 28478 6078 28530 6130
rect 29374 6078 29426 6130
rect 29598 6078 29650 6130
rect 33854 6078 33906 6130
rect 34190 6078 34242 6130
rect 38222 6078 38274 6130
rect 40238 6078 40290 6130
rect 41694 6078 41746 6130
rect 41806 6078 41858 6130
rect 5518 5966 5570 6018
rect 8878 5966 8930 6018
rect 11566 5966 11618 6018
rect 12350 5966 12402 6018
rect 15822 5966 15874 6018
rect 16830 5966 16882 6018
rect 19630 5966 19682 6018
rect 22430 5966 22482 6018
rect 28590 5966 28642 6018
rect 29934 5966 29986 6018
rect 31502 5966 31554 6018
rect 31838 5966 31890 6018
rect 32734 5966 32786 6018
rect 32846 5966 32898 6018
rect 33630 5966 33682 6018
rect 34078 5966 34130 6018
rect 35422 5966 35474 6018
rect 39566 5966 39618 6018
rect 40126 5966 40178 6018
rect 1934 5854 1986 5906
rect 9886 5854 9938 5906
rect 9998 5854 10050 5906
rect 10222 5854 10274 5906
rect 11006 5854 11058 5906
rect 17726 5854 17778 5906
rect 23214 5854 23266 5906
rect 24222 5854 24274 5906
rect 24670 5854 24722 5906
rect 25678 5854 25730 5906
rect 26238 5854 26290 5906
rect 26462 5854 26514 5906
rect 27470 5854 27522 5906
rect 27694 5854 27746 5906
rect 28030 5854 28082 5906
rect 29262 5854 29314 5906
rect 29822 5854 29874 5906
rect 30382 5854 30434 5906
rect 30494 5854 30546 5906
rect 30718 5854 30770 5906
rect 30942 5854 30994 5906
rect 32062 5854 32114 5906
rect 32510 5854 32562 5906
rect 34638 5854 34690 5906
rect 38110 5854 38162 5906
rect 38558 5910 38610 5962
rect 41582 5966 41634 6018
rect 39342 5854 39394 5906
rect 40462 5854 40514 5906
rect 2606 5742 2658 5794
rect 4734 5742 4786 5794
rect 6750 5742 6802 5794
rect 7646 5742 7698 5794
rect 10110 5742 10162 5794
rect 13470 5742 13522 5794
rect 14142 5742 14194 5794
rect 14814 5742 14866 5794
rect 18510 5742 18562 5794
rect 20302 5742 20354 5794
rect 24558 5742 24610 5794
rect 27806 5742 27858 5794
rect 31614 5742 31666 5794
rect 37550 5742 37602 5794
rect 14254 5630 14306 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 5854 5294 5906 5346
rect 12014 5294 12066 5346
rect 20302 5294 20354 5346
rect 33630 5294 33682 5346
rect 35982 5294 36034 5346
rect 36318 5294 36370 5346
rect 1822 5182 1874 5234
rect 2606 5182 2658 5234
rect 4958 5182 5010 5234
rect 6414 5182 6466 5234
rect 8430 5182 8482 5234
rect 10558 5182 10610 5234
rect 14254 5182 14306 5234
rect 14814 5182 14866 5234
rect 17614 5182 17666 5234
rect 19742 5182 19794 5234
rect 24670 5182 24722 5234
rect 26798 5182 26850 5234
rect 30718 5182 30770 5234
rect 32846 5182 32898 5234
rect 33406 5182 33458 5234
rect 33966 5182 34018 5234
rect 36766 5182 36818 5234
rect 37550 5182 37602 5234
rect 37886 5182 37938 5234
rect 38334 5182 38386 5234
rect 41358 5182 41410 5234
rect 2270 5070 2322 5122
rect 11230 5070 11282 5122
rect 12574 5070 12626 5122
rect 16830 5070 16882 5122
rect 20526 5070 20578 5122
rect 23438 5070 23490 5122
rect 23998 5070 24050 5122
rect 28478 5070 28530 5122
rect 29934 5070 29986 5122
rect 34974 5070 35026 5122
rect 39902 5070 39954 5122
rect 40686 5070 40738 5122
rect 2494 4958 2546 5010
rect 2718 4958 2770 5010
rect 3838 4958 3890 5010
rect 5742 4958 5794 5010
rect 7422 4958 7474 5010
rect 11902 4958 11954 5010
rect 12126 4958 12178 5010
rect 12350 4958 12402 5010
rect 15934 4958 15986 5010
rect 21870 4958 21922 5010
rect 22430 4958 22482 5010
rect 23102 4958 23154 5010
rect 27470 4958 27522 5010
rect 35086 4958 35138 5010
rect 35422 4958 35474 5010
rect 36094 4958 36146 5010
rect 39006 4958 39058 5010
rect 2830 4846 2882 4898
rect 13694 4846 13746 4898
rect 22094 4846 22146 4898
rect 22206 4846 22258 4898
rect 22318 4846 22370 4898
rect 23214 4846 23266 4898
rect 35310 4846 35362 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 6750 4510 6802 4562
rect 6974 4510 7026 4562
rect 9774 4510 9826 4562
rect 29038 4510 29090 4562
rect 32734 4510 32786 4562
rect 40014 4510 40066 4562
rect 40686 4510 40738 4562
rect 1822 4398 1874 4450
rect 6526 4398 6578 4450
rect 7646 4398 7698 4450
rect 9886 4398 9938 4450
rect 18062 4398 18114 4450
rect 21646 4398 21698 4450
rect 24782 4398 24834 4450
rect 26462 4398 26514 4450
rect 32846 4398 32898 4450
rect 33630 4398 33682 4450
rect 35422 4398 35474 4450
rect 40238 4398 40290 4450
rect 41582 4398 41634 4450
rect 2046 4286 2098 4338
rect 5966 4286 6018 4338
rect 10558 4286 10610 4338
rect 13918 4286 13970 4338
rect 14702 4286 14754 4338
rect 18174 4286 18226 4338
rect 18398 4286 18450 4338
rect 18622 4286 18674 4338
rect 22430 4286 22482 4338
rect 23998 4286 24050 4338
rect 25790 4286 25842 4338
rect 30830 4286 30882 4338
rect 31390 4286 31442 4338
rect 31614 4286 31666 4338
rect 31950 4286 32002 4338
rect 32510 4286 32562 4338
rect 33854 4286 33906 4338
rect 34638 4286 34690 4338
rect 39342 4286 39394 4338
rect 41806 4286 41858 4338
rect 3054 4174 3106 4226
rect 5182 4174 5234 4226
rect 8990 4174 9042 4226
rect 11230 4174 11282 4226
rect 13358 4174 13410 4226
rect 16830 4174 16882 4226
rect 19518 4174 19570 4226
rect 23102 4174 23154 4226
rect 28590 4174 28642 4226
rect 29710 4174 29762 4226
rect 37550 4174 37602 4226
rect 38222 4174 38274 4226
rect 7086 4062 7138 4114
rect 18734 4062 18786 4114
rect 24894 4062 24946 4114
rect 39902 4062 39954 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 4958 3726 5010 3778
rect 6862 3726 6914 3778
rect 10110 3726 10162 3778
rect 10334 3726 10386 3778
rect 10558 3726 10610 3778
rect 10670 3726 10722 3778
rect 14030 3726 14082 3778
rect 14254 3726 14306 3778
rect 14478 3726 14530 3778
rect 17726 3726 17778 3778
rect 23550 3726 23602 3778
rect 23886 3726 23938 3778
rect 41918 3726 41970 3778
rect 4174 3614 4226 3666
rect 4846 3614 4898 3666
rect 5854 3614 5906 3666
rect 6750 3614 6802 3666
rect 8878 3614 8930 3666
rect 12798 3614 12850 3666
rect 14590 3614 14642 3666
rect 15486 3614 15538 3666
rect 19182 3614 19234 3666
rect 21534 3614 21586 3666
rect 24446 3614 24498 3666
rect 27806 3614 27858 3666
rect 29934 3614 29986 3666
rect 33854 3614 33906 3666
rect 35646 3614 35698 3666
rect 40910 3614 40962 3666
rect 41582 3614 41634 3666
rect 5966 3502 6018 3554
rect 6190 3502 6242 3554
rect 17614 3502 17666 3554
rect 18286 3502 18338 3554
rect 18622 3502 18674 3554
rect 26350 3502 26402 3554
rect 27246 3502 27298 3554
rect 29486 3502 29538 3554
rect 32286 3502 32338 3554
rect 33182 3502 33234 3554
rect 34974 3502 35026 3554
rect 38334 3502 38386 3554
rect 40126 3502 40178 3554
rect 2270 3390 2322 3442
rect 7870 3390 7922 3442
rect 11678 3390 11730 3442
rect 13918 3390 13970 3442
rect 16606 3390 16658 3442
rect 20190 3390 20242 3442
rect 22542 3390 22594 3442
rect 23774 3390 23826 3442
rect 25454 3390 25506 3442
rect 31166 3390 31218 3442
rect 37214 3390 37266 3442
rect 39006 3390 39058 3442
rect 41694 3390 41746 3442
rect 6414 3278 6466 3330
rect 10222 3278 10274 3330
rect 17726 3278 17778 3330
rect 18510 3278 18562 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 15932 32340 15988 32350
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 2492 25508 2548 25518
rect 2492 25414 2548 25452
rect 1708 25396 1764 25406
rect 1484 25284 1540 25294
rect 1372 23716 1428 23726
rect 1148 23604 1204 23614
rect 1036 16772 1092 16782
rect 1036 3108 1092 16716
rect 1148 11396 1204 23548
rect 1148 11330 1204 11340
rect 1260 22372 1316 22382
rect 1260 6020 1316 22316
rect 1260 5954 1316 5964
rect 1372 5124 1428 23660
rect 1484 6580 1540 25228
rect 1484 6514 1540 6524
rect 1596 23828 1652 23838
rect 1372 5058 1428 5068
rect 1596 4900 1652 23772
rect 1708 19794 1764 25340
rect 13468 25396 13524 25406
rect 2940 25284 2996 25294
rect 2940 25190 2996 25228
rect 5068 25282 5124 25294
rect 5740 25284 5796 25294
rect 5068 25230 5070 25282
rect 5122 25230 5124 25282
rect 5068 24836 5124 25230
rect 4956 24780 5124 24836
rect 5628 25282 5796 25284
rect 5628 25230 5742 25282
rect 5794 25230 5796 25282
rect 5628 25228 5796 25230
rect 2268 24724 2324 24734
rect 1820 24610 1876 24622
rect 1820 24558 1822 24610
rect 1874 24558 1876 24610
rect 1820 23268 1876 24558
rect 1932 23716 1988 23726
rect 1932 23622 1988 23660
rect 2156 23380 2212 23390
rect 2156 23286 2212 23324
rect 1820 23212 1988 23268
rect 1820 23044 1876 23054
rect 1820 22950 1876 22988
rect 1820 22596 1876 22606
rect 1820 22482 1876 22540
rect 1820 22430 1822 22482
rect 1874 22430 1876 22482
rect 1820 22418 1876 22430
rect 1932 21252 1988 23212
rect 2268 22260 2324 24668
rect 2716 24612 2772 24622
rect 2716 24518 2772 24556
rect 3276 24610 3332 24622
rect 3276 24558 3278 24610
rect 3330 24558 3332 24610
rect 3276 23940 3332 24558
rect 4060 24610 4116 24622
rect 4060 24558 4062 24610
rect 4114 24558 4116 24610
rect 3276 23874 3332 23884
rect 3836 24500 3892 24510
rect 3724 23828 3780 23838
rect 3724 23734 3780 23772
rect 2380 23716 2436 23726
rect 2380 23714 2548 23716
rect 2380 23662 2382 23714
rect 2434 23662 2548 23714
rect 2380 23660 2548 23662
rect 2380 23650 2436 23660
rect 2268 22204 2436 22260
rect 2156 22148 2212 22158
rect 2156 22054 2212 22092
rect 1708 19742 1710 19794
rect 1762 19742 1764 19794
rect 1708 18340 1764 19742
rect 1820 21196 1988 21252
rect 2156 21474 2212 21486
rect 2156 21422 2158 21474
rect 2210 21422 2212 21474
rect 1820 19458 1876 21196
rect 1932 21026 1988 21038
rect 1932 20974 1934 21026
rect 1986 20974 1988 21026
rect 1932 20244 1988 20974
rect 2044 20692 2100 20702
rect 2044 20598 2100 20636
rect 1932 20242 2100 20244
rect 1932 20190 1934 20242
rect 1986 20190 2100 20242
rect 1932 20188 2100 20190
rect 1932 20178 1988 20188
rect 1820 19406 1822 19458
rect 1874 19406 1876 19458
rect 1820 19394 1876 19406
rect 1932 19460 1988 19470
rect 1932 19346 1988 19404
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1708 18274 1764 18284
rect 1820 18452 1876 18462
rect 1820 16996 1876 18396
rect 1932 17780 1988 19294
rect 2044 18116 2100 20188
rect 2156 19012 2212 21422
rect 2380 20914 2436 22204
rect 2492 21924 2548 23660
rect 2828 23714 2884 23726
rect 2828 23662 2830 23714
rect 2882 23662 2884 23714
rect 2716 23156 2772 23166
rect 2604 23044 2660 23054
rect 2604 22950 2660 22988
rect 2716 22482 2772 23100
rect 2716 22430 2718 22482
rect 2770 22430 2772 22482
rect 2716 22418 2772 22430
rect 2828 22036 2884 23662
rect 3276 23714 3332 23726
rect 3276 23662 3278 23714
rect 3330 23662 3332 23714
rect 3276 23604 3332 23662
rect 3276 23538 3332 23548
rect 3052 23380 3108 23390
rect 3052 22482 3108 23324
rect 3164 23042 3220 23054
rect 3164 22990 3166 23042
rect 3218 22990 3220 23042
rect 3164 22932 3220 22990
rect 3612 23044 3668 23054
rect 3612 23042 3780 23044
rect 3612 22990 3614 23042
rect 3666 22990 3780 23042
rect 3612 22988 3780 22990
rect 3612 22978 3668 22988
rect 3164 22866 3220 22876
rect 3052 22430 3054 22482
rect 3106 22430 3108 22482
rect 3052 22418 3108 22430
rect 3612 22146 3668 22158
rect 3612 22094 3614 22146
rect 3666 22094 3668 22146
rect 2828 21980 3220 22036
rect 2492 21868 2996 21924
rect 2492 21026 2548 21868
rect 2940 21810 2996 21868
rect 2940 21758 2942 21810
rect 2994 21758 2996 21810
rect 2940 21746 2996 21758
rect 2492 20974 2494 21026
rect 2546 20974 2548 21026
rect 2492 20962 2548 20974
rect 2604 21474 2660 21486
rect 2604 21422 2606 21474
rect 2658 21422 2660 21474
rect 2380 20862 2382 20914
rect 2434 20862 2436 20914
rect 2380 20244 2436 20862
rect 2604 20244 2660 21422
rect 2828 21362 2884 21374
rect 2828 21310 2830 21362
rect 2882 21310 2884 21362
rect 2828 20578 2884 21310
rect 2828 20526 2830 20578
rect 2882 20526 2884 20578
rect 2716 20244 2772 20254
rect 2604 20188 2716 20244
rect 2380 20178 2436 20188
rect 2716 20112 2772 20188
rect 2492 20020 2548 20030
rect 2268 19906 2324 19918
rect 2268 19854 2270 19906
rect 2322 19854 2324 19906
rect 2268 19794 2324 19854
rect 2268 19742 2270 19794
rect 2322 19742 2324 19794
rect 2268 19730 2324 19742
rect 2268 19124 2324 19134
rect 2268 19030 2324 19068
rect 2492 19124 2548 19964
rect 2828 20020 2884 20526
rect 2828 19954 2884 19964
rect 2940 20580 2996 20590
rect 2156 18946 2212 18956
rect 2156 18340 2212 18350
rect 2156 18246 2212 18284
rect 2380 18228 2436 18238
rect 2044 18060 2212 18116
rect 2044 17780 2100 17790
rect 1932 17778 2100 17780
rect 1932 17726 2046 17778
rect 2098 17726 2100 17778
rect 1932 17724 2100 17726
rect 2044 17714 2100 17724
rect 2044 17108 2100 17118
rect 1932 16996 1988 17006
rect 1820 16940 1932 16996
rect 1708 16884 1764 16894
rect 1932 16864 1988 16940
rect 1708 8372 1764 16828
rect 2044 16212 2100 17052
rect 1932 16156 2100 16212
rect 1820 16100 1876 16110
rect 1820 16006 1876 16044
rect 1932 15426 1988 16156
rect 2044 15540 2100 15550
rect 2156 15540 2212 18060
rect 2268 16882 2324 16894
rect 2268 16830 2270 16882
rect 2322 16830 2324 16882
rect 2268 16660 2324 16830
rect 2268 16594 2324 16604
rect 2380 16322 2436 18172
rect 2380 16270 2382 16322
rect 2434 16270 2436 16322
rect 2380 16258 2436 16270
rect 2268 16100 2324 16110
rect 2492 16100 2548 19068
rect 2828 19458 2884 19470
rect 2828 19406 2830 19458
rect 2882 19406 2884 19458
rect 2716 19012 2772 19022
rect 2716 18918 2772 18956
rect 2716 18338 2772 18350
rect 2716 18286 2718 18338
rect 2770 18286 2772 18338
rect 2716 17780 2772 18286
rect 2604 17668 2660 17678
rect 2604 17574 2660 17612
rect 2716 17332 2772 17724
rect 2828 17556 2884 19406
rect 2828 17490 2884 17500
rect 2716 17276 2884 17332
rect 2268 16098 2548 16100
rect 2268 16046 2270 16098
rect 2322 16046 2548 16098
rect 2268 16044 2548 16046
rect 2268 16034 2324 16044
rect 2044 15538 2212 15540
rect 2044 15486 2046 15538
rect 2098 15486 2212 15538
rect 2044 15484 2212 15486
rect 2044 15474 2100 15484
rect 1932 15374 1934 15426
rect 1986 15374 1988 15426
rect 1932 15316 1988 15374
rect 1932 15250 1988 15260
rect 2156 15148 2212 15484
rect 2268 15876 2324 15886
rect 2268 15538 2324 15820
rect 2268 15486 2270 15538
rect 2322 15486 2324 15538
rect 2268 15474 2324 15486
rect 2380 15874 2436 15886
rect 2380 15822 2382 15874
rect 2434 15822 2436 15874
rect 2380 15764 2436 15822
rect 2380 15316 2436 15708
rect 2044 15092 2212 15148
rect 2268 15260 2436 15316
rect 2044 14420 2100 15092
rect 2156 14644 2212 14654
rect 2156 14550 2212 14588
rect 2044 14364 2212 14420
rect 1932 13636 1988 13646
rect 1820 13580 1932 13636
rect 1820 12290 1876 13580
rect 1932 13542 1988 13580
rect 2044 13524 2100 13534
rect 2044 12962 2100 13468
rect 2044 12910 2046 12962
rect 2098 12910 2100 12962
rect 1932 12516 1988 12526
rect 1932 12402 1988 12460
rect 1932 12350 1934 12402
rect 1986 12350 1988 12402
rect 1932 12338 1988 12350
rect 1820 12238 1822 12290
rect 1874 12238 1876 12290
rect 1820 12226 1876 12238
rect 1820 11732 1876 11742
rect 1820 11506 1876 11676
rect 1820 11454 1822 11506
rect 1874 11454 1876 11506
rect 1820 11442 1876 11454
rect 1932 11060 1988 11070
rect 1932 10722 1988 11004
rect 1932 10670 1934 10722
rect 1986 10670 1988 10722
rect 1932 10658 1988 10670
rect 1820 9716 1876 9726
rect 2044 9716 2100 12910
rect 2156 12292 2212 14364
rect 2268 14196 2324 15260
rect 2492 15148 2548 16044
rect 2604 17108 2660 17118
rect 2604 15428 2660 17052
rect 2828 17106 2884 17276
rect 2828 17054 2830 17106
rect 2882 17054 2884 17106
rect 2828 17042 2884 17054
rect 2940 17108 2996 20524
rect 3164 20132 3220 21980
rect 3500 21476 3556 21486
rect 3500 21382 3556 21420
rect 3612 21362 3668 22094
rect 3612 21310 3614 21362
rect 3666 21310 3668 21362
rect 3612 21298 3668 21310
rect 3500 20692 3556 20702
rect 3500 20578 3556 20636
rect 3500 20526 3502 20578
rect 3554 20526 3556 20578
rect 3052 20130 3220 20132
rect 3052 20078 3166 20130
rect 3218 20078 3220 20130
rect 3052 20076 3220 20078
rect 3052 17892 3108 20076
rect 3164 20066 3220 20076
rect 3276 20244 3332 20254
rect 3164 19458 3220 19470
rect 3164 19406 3166 19458
rect 3218 19406 3220 19458
rect 3164 19346 3220 19406
rect 3164 19294 3166 19346
rect 3218 19294 3220 19346
rect 3164 19282 3220 19294
rect 3164 18340 3220 18350
rect 3164 18246 3220 18284
rect 3108 17836 3220 17892
rect 3052 17826 3108 17836
rect 3052 17444 3108 17454
rect 3052 17350 3108 17388
rect 3052 17108 3108 17118
rect 2940 17106 3108 17108
rect 2940 17054 3054 17106
rect 3106 17054 3108 17106
rect 2940 17052 3108 17054
rect 2716 16996 2772 17006
rect 2716 16902 2772 16940
rect 2828 15876 2884 15886
rect 2828 15538 2884 15820
rect 2828 15486 2830 15538
rect 2882 15486 2884 15538
rect 2716 15428 2772 15438
rect 2604 15426 2772 15428
rect 2604 15374 2718 15426
rect 2770 15374 2772 15426
rect 2604 15372 2772 15374
rect 2268 14130 2324 14140
rect 2380 15092 2548 15148
rect 2380 14530 2436 15092
rect 2380 14478 2382 14530
rect 2434 14478 2436 14530
rect 2268 12852 2324 12862
rect 2268 12758 2324 12796
rect 2156 12226 2212 12236
rect 2380 10164 2436 14478
rect 2492 12852 2548 12862
rect 2492 12290 2548 12796
rect 2604 12404 2660 12414
rect 2604 12310 2660 12348
rect 2492 12238 2494 12290
rect 2546 12238 2548 12290
rect 2492 11956 2548 12238
rect 2492 11890 2548 11900
rect 2604 12180 2660 12190
rect 2604 11732 2660 12124
rect 2380 10098 2436 10108
rect 2492 11676 2660 11732
rect 2156 9940 2212 9978
rect 2156 9874 2212 9884
rect 1820 9622 1876 9660
rect 1932 9714 2100 9716
rect 1932 9662 2046 9714
rect 2098 9662 2100 9714
rect 1932 9660 2100 9662
rect 1820 8932 1876 8942
rect 1932 8932 1988 9660
rect 2044 9650 2100 9660
rect 2156 9716 2212 9726
rect 2492 9716 2548 11676
rect 2716 10612 2772 15372
rect 2828 12740 2884 15486
rect 2940 15148 2996 17052
rect 3052 17042 3108 17052
rect 3164 17108 3220 17836
rect 3164 17042 3220 17052
rect 3276 16884 3332 20188
rect 3500 20132 3556 20526
rect 3724 20356 3780 22988
rect 3836 21812 3892 24444
rect 3948 23042 4004 23054
rect 3948 22990 3950 23042
rect 4002 22990 4004 23042
rect 3948 22594 4004 22990
rect 3948 22542 3950 22594
rect 4002 22542 4004 22594
rect 3948 22530 4004 22542
rect 4060 22372 4116 24558
rect 4508 24610 4564 24622
rect 4508 24558 4510 24610
rect 4562 24558 4564 24610
rect 4508 24500 4564 24558
rect 4956 24612 5012 24780
rect 4508 24444 4900 24500
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4172 23714 4228 23726
rect 4172 23662 4174 23714
rect 4226 23662 4228 23714
rect 4172 23492 4228 23662
rect 4620 23716 4676 23726
rect 4620 23622 4676 23660
rect 4396 23492 4452 23502
rect 4172 23436 4396 23492
rect 4396 23044 4452 23436
rect 4284 23042 4452 23044
rect 4284 22990 4398 23042
rect 4450 22990 4452 23042
rect 4284 22988 4452 22990
rect 4284 22484 4340 22988
rect 4396 22978 4452 22988
rect 4844 23044 4900 24444
rect 4956 23716 5012 24556
rect 5068 24612 5124 24622
rect 5516 24612 5572 24622
rect 5068 24610 5348 24612
rect 5068 24558 5070 24610
rect 5122 24558 5348 24610
rect 5068 24556 5348 24558
rect 5068 24546 5124 24556
rect 4956 23622 5012 23660
rect 4844 23042 5012 23044
rect 4844 22990 4846 23042
rect 4898 22990 5012 23042
rect 4844 22988 5012 22990
rect 4844 22978 4900 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4956 22594 5012 22988
rect 4956 22542 4958 22594
rect 5010 22542 5012 22594
rect 4396 22484 4452 22494
rect 4284 22482 4452 22484
rect 4284 22430 4398 22482
rect 4450 22430 4452 22482
rect 4284 22428 4452 22430
rect 4396 22418 4452 22428
rect 4844 22484 4900 22494
rect 4060 22306 4116 22316
rect 3836 21746 3892 21756
rect 4060 22146 4116 22158
rect 4060 22094 4062 22146
rect 4114 22094 4116 22146
rect 4060 21812 4116 22094
rect 3836 21588 3892 21598
rect 3836 21494 3892 21532
rect 3948 20692 4004 20702
rect 3948 20578 4004 20636
rect 3948 20526 3950 20578
rect 4002 20526 4004 20578
rect 3948 20468 4004 20526
rect 3948 20402 4004 20412
rect 3724 20290 3780 20300
rect 4060 20244 4116 21756
rect 4732 21812 4788 21822
rect 4732 21718 4788 21756
rect 4284 21700 4340 21710
rect 4284 21606 4340 21644
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4732 20804 4788 20814
rect 4620 20580 4676 20590
rect 4620 20486 4676 20524
rect 3948 20188 4060 20244
rect 3500 20076 3892 20132
rect 3500 19460 3556 19470
rect 3500 18674 3556 19404
rect 3500 18622 3502 18674
rect 3554 18622 3556 18674
rect 3388 18452 3444 18462
rect 3388 17778 3444 18396
rect 3388 17726 3390 17778
rect 3442 17726 3444 17778
rect 3388 17714 3444 17726
rect 3500 17332 3556 18622
rect 3500 17266 3556 17276
rect 3612 19012 3668 19022
rect 3612 18226 3668 18956
rect 3836 18340 3892 20076
rect 3948 19348 4004 20188
rect 4060 20178 4116 20188
rect 4284 20244 4340 20254
rect 4060 19906 4116 19918
rect 4060 19854 4062 19906
rect 4114 19854 4116 19906
rect 4060 19796 4116 19854
rect 4116 19740 4228 19796
rect 4060 19730 4116 19740
rect 4060 19348 4116 19358
rect 3948 19346 4116 19348
rect 3948 19294 4062 19346
rect 4114 19294 4116 19346
rect 3948 19292 4116 19294
rect 4060 19282 4116 19292
rect 3948 18340 4004 18350
rect 3836 18338 4004 18340
rect 3836 18286 3950 18338
rect 4002 18286 4004 18338
rect 3836 18284 4004 18286
rect 3612 18174 3614 18226
rect 3666 18174 3668 18226
rect 3052 16828 3332 16884
rect 3052 16100 3108 16828
rect 3500 16212 3556 16222
rect 3052 16098 3332 16100
rect 3052 16046 3054 16098
rect 3106 16046 3332 16098
rect 3052 16044 3332 16046
rect 3052 16034 3108 16044
rect 3164 15876 3220 15886
rect 3164 15782 3220 15820
rect 3052 15540 3108 15550
rect 3052 15446 3108 15484
rect 2940 15092 3108 15148
rect 2940 14306 2996 14318
rect 2940 14254 2942 14306
rect 2994 14254 2996 14306
rect 2940 12964 2996 14254
rect 3052 13188 3108 15092
rect 3052 13122 3108 13132
rect 2940 12898 2996 12908
rect 3164 12964 3220 12974
rect 3276 12964 3332 16044
rect 3388 15876 3444 15886
rect 3388 15782 3444 15820
rect 3500 15426 3556 16156
rect 3612 15764 3668 18174
rect 3948 18116 4004 18284
rect 3948 18050 4004 18060
rect 4060 17892 4116 17902
rect 4172 17892 4228 19740
rect 4060 17890 4228 17892
rect 4060 17838 4062 17890
rect 4114 17838 4228 17890
rect 4060 17836 4228 17838
rect 4284 18340 4340 20188
rect 4732 20242 4788 20748
rect 4732 20190 4734 20242
rect 4786 20190 4788 20242
rect 4732 20178 4788 20190
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19010 4676 19022
rect 4620 18958 4622 19010
rect 4674 18958 4676 19010
rect 4620 18900 4676 18958
rect 4620 18834 4676 18844
rect 4844 18674 4900 22428
rect 4956 20916 5012 22542
rect 4956 20850 5012 20860
rect 5068 20578 5124 20590
rect 5068 20526 5070 20578
rect 5122 20526 5124 20578
rect 5068 19908 5124 20526
rect 5068 19842 5124 19852
rect 5180 19906 5236 19918
rect 5180 19854 5182 19906
rect 5234 19854 5236 19906
rect 5180 19460 5236 19854
rect 5292 19572 5348 24556
rect 5404 24610 5572 24612
rect 5404 24558 5518 24610
rect 5570 24558 5572 24610
rect 5404 24556 5572 24558
rect 5404 23044 5460 24556
rect 5516 24546 5572 24556
rect 5628 23380 5684 25228
rect 5740 25218 5796 25228
rect 6188 25282 6244 25294
rect 6188 25230 6190 25282
rect 6242 25230 6244 25282
rect 5964 24612 6020 24622
rect 5964 24610 6132 24612
rect 5964 24558 5966 24610
rect 6018 24558 6132 24610
rect 5964 24556 6132 24558
rect 5964 24546 6020 24556
rect 5964 23940 6020 23950
rect 5740 23828 5796 23838
rect 5740 23734 5796 23772
rect 5740 23380 5796 23390
rect 5628 23324 5740 23380
rect 5404 22978 5460 22988
rect 5516 23042 5572 23054
rect 5516 22990 5518 23042
rect 5570 22990 5572 23042
rect 5516 22148 5572 22990
rect 5740 22260 5796 23324
rect 5740 22194 5796 22204
rect 5404 21588 5460 21598
rect 5404 21494 5460 21532
rect 5516 20804 5572 22092
rect 5740 21812 5796 21822
rect 5740 21718 5796 21756
rect 5516 20738 5572 20748
rect 5628 21476 5684 21486
rect 5628 20914 5684 21420
rect 5628 20862 5630 20914
rect 5682 20862 5684 20914
rect 5628 20132 5684 20862
rect 5964 20468 6020 23884
rect 6076 22484 6132 24556
rect 6188 24052 6244 25230
rect 6972 25282 7028 25294
rect 6972 25230 6974 25282
rect 7026 25230 7028 25282
rect 6860 24724 6916 24734
rect 6860 24630 6916 24668
rect 6412 24610 6468 24622
rect 6412 24558 6414 24610
rect 6466 24558 6468 24610
rect 6412 24164 6468 24558
rect 6412 24098 6468 24108
rect 6188 23986 6244 23996
rect 6300 23714 6356 23726
rect 6300 23662 6302 23714
rect 6354 23662 6356 23714
rect 6300 23156 6356 23662
rect 6860 23714 6916 23726
rect 6860 23662 6862 23714
rect 6914 23662 6916 23714
rect 6860 23604 6916 23662
rect 6860 23538 6916 23548
rect 6300 23090 6356 23100
rect 6860 23156 6916 23166
rect 6972 23156 7028 25230
rect 7420 25284 7476 25294
rect 7420 25282 7588 25284
rect 7420 25230 7422 25282
rect 7474 25230 7588 25282
rect 7420 25228 7588 25230
rect 7420 25218 7476 25228
rect 6916 23100 7028 23156
rect 7308 24610 7364 24622
rect 7308 24558 7310 24610
rect 7362 24558 7364 24610
rect 6860 23090 6916 23100
rect 6188 23042 6244 23054
rect 6188 22990 6190 23042
rect 6242 22990 6244 23042
rect 6188 22708 6244 22990
rect 6188 22642 6244 22652
rect 6412 23044 6468 23054
rect 6076 22418 6132 22428
rect 6300 22260 6356 22270
rect 5964 20402 6020 20412
rect 6076 22146 6132 22158
rect 6076 22094 6078 22146
rect 6130 22094 6132 22146
rect 6076 21812 6132 22094
rect 6188 21812 6244 21822
rect 6076 21810 6244 21812
rect 6076 21758 6190 21810
rect 6242 21758 6244 21810
rect 6076 21756 6244 21758
rect 6076 20244 6132 21756
rect 6188 21746 6244 21756
rect 6300 21588 6356 22204
rect 6076 20178 6132 20188
rect 6188 21532 6356 21588
rect 6412 22146 6468 22988
rect 6412 22094 6414 22146
rect 6466 22094 6468 22146
rect 5628 20066 5684 20076
rect 5964 19908 6020 19918
rect 6188 19908 6244 21532
rect 6300 20580 6356 20590
rect 6300 20486 6356 20524
rect 5964 19906 6244 19908
rect 5964 19854 5966 19906
rect 6018 19854 6244 19906
rect 5964 19852 6244 19854
rect 6412 19908 6468 22094
rect 6524 23042 6580 23054
rect 7084 23044 7140 23054
rect 6524 22990 6526 23042
rect 6578 22990 6580 23042
rect 6524 22932 6580 22990
rect 6524 21924 6580 22876
rect 6972 23042 7140 23044
rect 6972 22990 7086 23042
rect 7138 22990 7140 23042
rect 6972 22988 7140 22990
rect 6524 21858 6580 21868
rect 6860 22146 6916 22158
rect 6860 22094 6862 22146
rect 6914 22094 6916 22146
rect 6860 21924 6916 22094
rect 6860 21858 6916 21868
rect 6748 21474 6804 21486
rect 6748 21422 6750 21474
rect 6802 21422 6804 21474
rect 5964 19684 6020 19852
rect 6412 19842 6468 19852
rect 6524 21364 6580 21374
rect 5292 19516 5796 19572
rect 5180 19394 5236 19404
rect 5740 19458 5796 19516
rect 5740 19406 5742 19458
rect 5794 19406 5796 19458
rect 5740 19346 5796 19406
rect 5740 19294 5742 19346
rect 5794 19294 5796 19346
rect 5068 19012 5124 19022
rect 4844 18622 4846 18674
rect 4898 18622 4900 18674
rect 4284 17892 4340 18284
rect 4396 18338 4452 18350
rect 4396 18286 4398 18338
rect 4450 18286 4452 18338
rect 4396 18226 4452 18286
rect 4844 18340 4900 18622
rect 4956 19010 5124 19012
rect 4956 18958 5070 19010
rect 5122 18958 5124 19010
rect 4956 18956 5124 18958
rect 4956 18564 5012 18956
rect 5068 18946 5124 18956
rect 4956 18498 5012 18508
rect 5068 18788 5124 18798
rect 4844 18274 4900 18284
rect 4396 18174 4398 18226
rect 4450 18174 4452 18226
rect 4396 18162 4452 18174
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 5068 18004 5124 18732
rect 5292 18340 5348 18350
rect 5292 18246 5348 18284
rect 4476 17994 4740 18004
rect 4844 17948 5124 18004
rect 4284 17836 4564 17892
rect 4060 17826 4116 17836
rect 3948 17554 4004 17566
rect 3948 17502 3950 17554
rect 4002 17502 4004 17554
rect 3724 16996 3780 17006
rect 3724 16100 3780 16940
rect 3836 16884 3892 16894
rect 3836 16790 3892 16828
rect 3948 16324 4004 17502
rect 3948 16258 4004 16268
rect 4172 16212 4228 17836
rect 4396 17668 4452 17678
rect 4396 17220 4452 17612
rect 4396 16994 4452 17164
rect 4396 16942 4398 16994
rect 4450 16942 4452 16994
rect 4396 16930 4452 16942
rect 4508 17106 4564 17836
rect 4844 17890 4900 17948
rect 4844 17838 4846 17890
rect 4898 17838 4900 17890
rect 4844 17826 4900 17838
rect 5628 17668 5684 17678
rect 5628 17574 5684 17612
rect 4956 17554 5012 17566
rect 4956 17502 4958 17554
rect 5010 17502 5012 17554
rect 4844 17444 4900 17454
rect 4844 17350 4900 17388
rect 4508 17054 4510 17106
rect 4562 17054 4564 17106
rect 4508 16660 4564 17054
rect 4956 17108 5012 17502
rect 4956 17042 5012 17052
rect 5292 17444 5348 17454
rect 5292 17106 5348 17388
rect 5292 17054 5294 17106
rect 5346 17054 5348 17106
rect 5292 17042 5348 17054
rect 5404 17332 5460 17342
rect 5068 16996 5124 17006
rect 5068 16902 5124 16940
rect 5404 16994 5460 17276
rect 5404 16942 5406 16994
rect 5458 16942 5460 16994
rect 5404 16930 5460 16942
rect 4732 16884 4788 16894
rect 4732 16882 5012 16884
rect 4732 16830 4734 16882
rect 4786 16830 5012 16882
rect 4732 16828 5012 16830
rect 4732 16818 4788 16828
rect 4284 16604 4564 16660
rect 4284 16324 4340 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16436 4900 16446
rect 4732 16324 4788 16334
rect 4284 16268 4564 16324
rect 4172 16156 4452 16212
rect 3836 16100 3892 16110
rect 3724 16098 4340 16100
rect 3724 16046 3838 16098
rect 3890 16046 4340 16098
rect 3724 16044 4340 16046
rect 3836 16034 3892 16044
rect 3948 15930 4004 15942
rect 3836 15876 3892 15886
rect 3948 15878 3950 15930
rect 4002 15878 4004 15930
rect 3948 15876 4004 15878
rect 3892 15820 4004 15876
rect 4172 15874 4228 15886
rect 4172 15822 4174 15874
rect 4226 15822 4228 15874
rect 3836 15810 3892 15820
rect 3612 15698 3668 15708
rect 4060 15764 4116 15774
rect 3500 15374 3502 15426
rect 3554 15374 3556 15426
rect 3500 15362 3556 15374
rect 3612 15428 3668 15438
rect 3612 15426 3780 15428
rect 3612 15374 3614 15426
rect 3666 15374 3780 15426
rect 3612 15372 3780 15374
rect 3612 15362 3668 15372
rect 3500 14420 3556 14430
rect 3500 14326 3556 14364
rect 3612 14308 3668 14318
rect 3164 12962 3332 12964
rect 3164 12910 3166 12962
rect 3218 12910 3332 12962
rect 3164 12908 3332 12910
rect 3164 12898 3220 12908
rect 3276 12852 3332 12908
rect 3052 12740 3108 12750
rect 2828 12684 2996 12740
rect 2828 12180 2884 12190
rect 2828 12086 2884 12124
rect 1820 8930 2100 8932
rect 1820 8878 1822 8930
rect 1874 8878 2100 8930
rect 1820 8876 2100 8878
rect 1820 8866 1876 8876
rect 1932 8484 1988 8494
rect 1932 8390 1988 8428
rect 1820 8372 1876 8382
rect 1708 8370 1876 8372
rect 1708 8318 1822 8370
rect 1874 8318 1876 8370
rect 1708 8316 1876 8318
rect 1820 8306 1876 8316
rect 2044 8260 2100 8876
rect 2044 8194 2100 8204
rect 2156 8596 2212 9660
rect 1596 4834 1652 4844
rect 1708 8036 1764 8046
rect 2156 8036 2212 8540
rect 2380 9660 2548 9716
rect 2604 10556 2772 10612
rect 1708 4452 1764 7980
rect 1820 7980 2212 8036
rect 2268 8148 2324 8158
rect 1820 7362 1876 7980
rect 2044 7588 2100 7598
rect 1820 7310 1822 7362
rect 1874 7310 1876 7362
rect 1820 5684 1876 7310
rect 1932 7476 1988 7486
rect 1932 5906 1988 7420
rect 2044 6466 2100 7532
rect 2044 6414 2046 6466
rect 2098 6414 2100 6466
rect 2044 6402 2100 6414
rect 2156 6578 2212 6590
rect 2156 6526 2158 6578
rect 2210 6526 2212 6578
rect 1932 5854 1934 5906
rect 1986 5854 1988 5906
rect 1932 5842 1988 5854
rect 1820 5628 2100 5684
rect 1820 5236 1876 5246
rect 1820 5142 1876 5180
rect 1820 4452 1876 4462
rect 1708 4450 1876 4452
rect 1708 4398 1822 4450
rect 1874 4398 1876 4450
rect 1708 4396 1876 4398
rect 1820 4386 1876 4396
rect 2044 4338 2100 5628
rect 2156 4564 2212 6526
rect 2268 5122 2324 8092
rect 2380 8036 2436 9660
rect 2492 8260 2548 8270
rect 2604 8260 2660 10556
rect 2716 9940 2772 9950
rect 2716 9846 2772 9884
rect 2940 9828 2996 12684
rect 3052 12738 3220 12740
rect 3052 12686 3054 12738
rect 3106 12686 3220 12738
rect 3052 12684 3220 12686
rect 3052 12674 3108 12684
rect 3164 12180 3220 12684
rect 3164 12114 3220 12124
rect 3276 11732 3332 12796
rect 3388 12964 3444 12974
rect 3388 11788 3444 12908
rect 3500 12178 3556 12190
rect 3500 12126 3502 12178
rect 3554 12126 3556 12178
rect 3500 11956 3556 12126
rect 3500 11890 3556 11900
rect 3388 11732 3556 11788
rect 3276 11666 3332 11676
rect 3388 11508 3444 11518
rect 3164 11284 3220 11294
rect 2828 9772 2996 9828
rect 3052 9938 3108 9950
rect 3052 9886 3054 9938
rect 3106 9886 3108 9938
rect 3052 9828 3108 9886
rect 2492 8258 2660 8260
rect 2492 8206 2494 8258
rect 2546 8206 2660 8258
rect 2492 8204 2660 8206
rect 2716 8260 2772 8270
rect 2828 8260 2884 9772
rect 3052 9762 3108 9772
rect 2940 9602 2996 9614
rect 2940 9550 2942 9602
rect 2994 9550 2996 9602
rect 2940 8484 2996 9550
rect 2940 8418 2996 8428
rect 3052 8372 3108 8382
rect 3052 8278 3108 8316
rect 2716 8258 2884 8260
rect 2716 8206 2718 8258
rect 2770 8206 2884 8258
rect 2716 8204 2884 8206
rect 2492 8194 2548 8204
rect 2716 8194 2772 8204
rect 2380 7970 2436 7980
rect 2828 7812 2884 8204
rect 2940 8148 2996 8158
rect 3164 8148 3220 11228
rect 3276 10500 3332 10510
rect 3388 10500 3444 11452
rect 3276 10498 3444 10500
rect 3276 10446 3278 10498
rect 3330 10446 3444 10498
rect 3276 10444 3444 10446
rect 3276 10434 3332 10444
rect 3500 10276 3556 11732
rect 3612 10612 3668 14252
rect 3724 13076 3780 15372
rect 3836 15316 3892 15326
rect 3836 15314 4004 15316
rect 3836 15262 3838 15314
rect 3890 15262 4004 15314
rect 3836 15260 4004 15262
rect 3836 15250 3892 15260
rect 3948 15204 4004 15260
rect 3836 14756 3892 14766
rect 3836 14530 3892 14700
rect 3836 14478 3838 14530
rect 3890 14478 3892 14530
rect 3836 14466 3892 14478
rect 3948 13972 4004 15148
rect 3836 13916 4004 13972
rect 3836 13300 3892 13916
rect 4060 13860 4116 15708
rect 4172 15428 4228 15822
rect 4172 15362 4228 15372
rect 4284 15426 4340 16044
rect 4396 15538 4452 16156
rect 4508 15764 4564 16268
rect 4732 16210 4788 16268
rect 4732 16158 4734 16210
rect 4786 16158 4788 16210
rect 4732 16146 4788 16158
rect 4620 15986 4676 15998
rect 4620 15934 4622 15986
rect 4674 15934 4676 15986
rect 4620 15876 4676 15934
rect 4844 15986 4900 16380
rect 4844 15934 4846 15986
rect 4898 15934 4900 15986
rect 4844 15922 4900 15934
rect 4620 15810 4676 15820
rect 4508 15698 4564 15708
rect 4396 15486 4398 15538
rect 4450 15486 4452 15538
rect 4396 15474 4452 15486
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15362 4340 15374
rect 4620 15316 4676 15326
rect 4620 15222 4676 15260
rect 4844 15092 4900 15102
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4284 14418 4340 14430
rect 4284 14366 4286 14418
rect 4338 14366 4340 14418
rect 4284 14196 4340 14366
rect 4396 14308 4452 14318
rect 4396 14214 4452 14252
rect 4284 14130 4340 14140
rect 3836 13234 3892 13244
rect 3948 13804 4116 13860
rect 3724 13010 3780 13020
rect 3948 13074 4004 13804
rect 4844 13748 4900 15036
rect 4956 13972 5012 16828
rect 5740 16548 5796 19294
rect 5964 18452 6020 19628
rect 6188 19458 6244 19470
rect 6188 19406 6190 19458
rect 6242 19406 6244 19458
rect 6188 18564 6244 19406
rect 6300 19012 6356 19022
rect 6300 19010 6468 19012
rect 6300 18958 6302 19010
rect 6354 18958 6468 19010
rect 6300 18956 6468 18958
rect 6300 18946 6356 18956
rect 6300 18564 6356 18574
rect 6188 18562 6356 18564
rect 6188 18510 6302 18562
rect 6354 18510 6356 18562
rect 6188 18508 6356 18510
rect 6300 18498 6356 18508
rect 6412 18564 6468 18956
rect 6524 18788 6580 21308
rect 6748 21140 6804 21422
rect 6748 21074 6804 21084
rect 6636 20804 6692 20814
rect 6636 20578 6692 20748
rect 6972 20580 7028 22988
rect 7084 22978 7140 22988
rect 7196 22036 7252 22046
rect 7084 21476 7140 21486
rect 7196 21476 7252 21980
rect 7084 21474 7252 21476
rect 7084 21422 7086 21474
rect 7138 21422 7252 21474
rect 7084 21420 7252 21422
rect 7084 21410 7140 21420
rect 7084 20916 7140 20926
rect 7084 20822 7140 20860
rect 6636 20526 6638 20578
rect 6690 20526 6692 20578
rect 6636 19236 6692 20526
rect 6636 19170 6692 19180
rect 6748 20524 7028 20580
rect 6748 20130 6804 20524
rect 7196 20244 7252 21420
rect 6748 20078 6750 20130
rect 6802 20078 6804 20130
rect 6524 18722 6580 18732
rect 6636 19010 6692 19022
rect 6636 18958 6638 19010
rect 6690 18958 6692 19010
rect 6636 18676 6692 18958
rect 6636 18610 6692 18620
rect 6412 18498 6468 18508
rect 5964 18386 6020 18396
rect 6524 18452 6580 18462
rect 5852 18338 5908 18350
rect 5852 18286 5854 18338
rect 5906 18286 5908 18338
rect 5852 18004 5908 18286
rect 6412 18340 6468 18350
rect 6076 18228 6132 18238
rect 6076 18226 6244 18228
rect 6076 18174 6078 18226
rect 6130 18174 6244 18226
rect 6076 18172 6244 18174
rect 6076 18162 6132 18172
rect 5852 17938 5908 17948
rect 6188 17666 6244 18172
rect 6300 17892 6356 17902
rect 6300 17798 6356 17836
rect 6188 17614 6190 17666
rect 6242 17614 6244 17666
rect 6188 17602 6244 17614
rect 6076 17556 6132 17566
rect 5628 16492 5796 16548
rect 5852 17444 5908 17454
rect 5068 15988 5124 15998
rect 5068 15426 5124 15932
rect 5516 15988 5572 15998
rect 5180 15876 5236 15886
rect 5180 15538 5236 15820
rect 5180 15486 5182 15538
rect 5234 15486 5236 15538
rect 5180 15474 5236 15486
rect 5404 15540 5460 15550
rect 5404 15446 5460 15484
rect 5068 15374 5070 15426
rect 5122 15374 5124 15426
rect 5068 15362 5124 15374
rect 4956 13906 5012 13916
rect 5404 14756 5460 14766
rect 4060 13636 4116 13646
rect 4844 13616 4900 13692
rect 5180 13748 5236 13758
rect 4060 13542 4116 13580
rect 4844 13524 4900 13534
rect 4476 13356 4740 13366
rect 4060 13300 4116 13310
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4060 13188 4116 13244
rect 4620 13188 4676 13198
rect 4844 13188 4900 13468
rect 4060 13132 4564 13188
rect 3948 13022 3950 13074
rect 4002 13022 4004 13074
rect 3836 12738 3892 12750
rect 3836 12686 3838 12738
rect 3890 12686 3892 12738
rect 3724 12628 3780 12638
rect 3724 12402 3780 12572
rect 3724 12350 3726 12402
rect 3778 12350 3780 12402
rect 3724 12338 3780 12350
rect 3836 12404 3892 12686
rect 3948 12740 4004 13022
rect 4060 12852 4116 12862
rect 4396 12852 4452 12862
rect 4060 12850 4228 12852
rect 4060 12798 4062 12850
rect 4114 12798 4228 12850
rect 4060 12796 4228 12798
rect 4060 12786 4116 12796
rect 3948 12674 4004 12684
rect 3836 12338 3892 12348
rect 3948 12292 4004 12302
rect 3948 12198 4004 12236
rect 4172 12292 4228 12796
rect 4172 12226 4228 12236
rect 3724 12180 3780 12190
rect 3780 12124 3892 12180
rect 3724 12048 3780 12124
rect 3612 10546 3668 10556
rect 3724 11844 3780 11854
rect 3724 10500 3780 11788
rect 3836 10836 3892 12124
rect 4284 12068 4340 12078
rect 4396 12068 4452 12796
rect 4508 12290 4564 13132
rect 4620 13186 4900 13188
rect 4620 13134 4622 13186
rect 4674 13134 4900 13186
rect 4620 13132 4900 13134
rect 4620 13122 4676 13132
rect 5180 13076 5236 13692
rect 5404 13524 5460 14700
rect 5516 13746 5572 15932
rect 5516 13694 5518 13746
rect 5570 13694 5572 13746
rect 5516 13682 5572 13694
rect 5628 13748 5684 16492
rect 5740 16324 5796 16334
rect 5740 16230 5796 16268
rect 5852 16100 5908 17388
rect 6076 17108 6132 17500
rect 6300 17556 6356 17566
rect 6412 17556 6468 18284
rect 6524 17892 6580 18396
rect 6636 18450 6692 18462
rect 6636 18398 6638 18450
rect 6690 18398 6692 18450
rect 6636 18116 6692 18398
rect 6636 18050 6692 18060
rect 6524 17836 6692 17892
rect 6300 17554 6580 17556
rect 6300 17502 6302 17554
rect 6354 17502 6580 17554
rect 6300 17500 6580 17502
rect 6300 17490 6356 17500
rect 6188 17108 6244 17118
rect 6076 17106 6244 17108
rect 6076 17054 6190 17106
rect 6242 17054 6244 17106
rect 6076 17052 6244 17054
rect 6188 17042 6244 17052
rect 6412 16994 6468 17006
rect 6412 16942 6414 16994
rect 6466 16942 6468 16994
rect 5740 16044 5908 16100
rect 5964 16884 6020 16894
rect 5740 14756 5796 16044
rect 5964 15986 6020 16828
rect 6412 16772 6468 16942
rect 6524 16996 6580 17500
rect 6524 16864 6580 16940
rect 6412 16706 6468 16716
rect 6076 16324 6132 16334
rect 6076 16230 6132 16268
rect 5964 15934 5966 15986
rect 6018 15934 6020 15986
rect 5964 15922 6020 15934
rect 6524 16098 6580 16110
rect 6524 16046 6526 16098
rect 6578 16046 6580 16098
rect 5852 15428 5908 15438
rect 5852 15334 5908 15372
rect 6300 15428 6356 15438
rect 6300 15334 6356 15372
rect 6076 15314 6132 15326
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 6076 14980 6132 15262
rect 6076 14914 6132 14924
rect 6412 15314 6468 15326
rect 6412 15262 6414 15314
rect 6466 15262 6468 15314
rect 5740 14690 5796 14700
rect 6076 14532 6132 14542
rect 5740 14530 6132 14532
rect 5740 14478 6078 14530
rect 6130 14478 6132 14530
rect 5740 14476 6132 14478
rect 5740 14084 5796 14476
rect 6076 14466 6132 14476
rect 5852 14308 5908 14318
rect 5852 14214 5908 14252
rect 5964 14306 6020 14318
rect 5964 14254 5966 14306
rect 6018 14254 6020 14306
rect 5740 14028 5908 14084
rect 5628 13682 5684 13692
rect 5740 13634 5796 13646
rect 5740 13582 5742 13634
rect 5794 13582 5796 13634
rect 5404 13468 5684 13524
rect 4956 13020 5236 13076
rect 4844 12964 4900 12974
rect 4620 12908 4844 12964
rect 4620 12402 4676 12908
rect 4844 12898 4900 12908
rect 4620 12350 4622 12402
rect 4674 12350 4676 12402
rect 4620 12338 4676 12350
rect 4732 12738 4788 12750
rect 4732 12686 4734 12738
rect 4786 12686 4788 12738
rect 4508 12238 4510 12290
rect 4562 12238 4564 12290
rect 4508 12226 4564 12238
rect 4732 12292 4788 12686
rect 4732 12226 4788 12236
rect 4844 12738 4900 12750
rect 4844 12686 4846 12738
rect 4898 12686 4900 12738
rect 4844 12068 4900 12686
rect 4396 12012 4900 12068
rect 4284 11620 4340 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11732 4900 12012
rect 4844 11666 4900 11676
rect 4284 11564 4676 11620
rect 3948 11284 4004 11294
rect 3948 11282 4340 11284
rect 3948 11230 3950 11282
rect 4002 11230 4340 11282
rect 3948 11228 4340 11230
rect 3948 11218 4004 11228
rect 4172 10836 4228 10846
rect 3836 10834 4228 10836
rect 3836 10782 4174 10834
rect 4226 10782 4228 10834
rect 3836 10780 4228 10782
rect 4172 10770 4228 10780
rect 4284 10834 4340 11228
rect 4284 10782 4286 10834
rect 4338 10782 4340 10834
rect 4284 10770 4340 10782
rect 4396 10948 4452 10958
rect 4396 10834 4452 10892
rect 4396 10782 4398 10834
rect 4450 10782 4452 10834
rect 4396 10770 4452 10782
rect 4508 10836 4564 10846
rect 4508 10742 4564 10780
rect 3948 10610 4004 10622
rect 3948 10558 3950 10610
rect 4002 10558 4004 10610
rect 3724 10444 3892 10500
rect 3612 10276 3668 10286
rect 3500 10220 3612 10276
rect 2940 8146 3220 8148
rect 2940 8094 2942 8146
rect 2994 8094 3220 8146
rect 2940 8092 3220 8094
rect 3276 10052 3332 10062
rect 3276 9268 3332 9996
rect 3612 9716 3668 10220
rect 3836 9826 3892 10444
rect 3948 10276 4004 10558
rect 4172 10612 4228 10622
rect 4620 10612 4676 11564
rect 4956 11508 5012 13020
rect 5404 12964 5460 12974
rect 4732 11452 5012 11508
rect 5068 12628 5124 12638
rect 4732 11394 4788 11452
rect 4732 11342 4734 11394
rect 4786 11342 4788 11394
rect 4732 11330 4788 11342
rect 5068 11284 5124 12572
rect 5180 12404 5236 12414
rect 5180 12290 5236 12348
rect 5180 12238 5182 12290
rect 5234 12238 5236 12290
rect 5180 12226 5236 12238
rect 5404 12402 5460 12908
rect 5404 12350 5406 12402
rect 5458 12350 5460 12402
rect 5404 11788 5460 12350
rect 5628 12290 5684 13468
rect 5740 12962 5796 13582
rect 5740 12910 5742 12962
rect 5794 12910 5796 12962
rect 5740 12898 5796 12910
rect 5628 12238 5630 12290
rect 5682 12238 5684 12290
rect 5404 11732 5572 11788
rect 3948 10210 4004 10220
rect 4060 10388 4116 10398
rect 3836 9774 3838 9826
rect 3890 9774 3892 9826
rect 3836 9762 3892 9774
rect 4060 9826 4116 10332
rect 4172 9940 4228 10556
rect 4172 9874 4228 9884
rect 4284 10556 4676 10612
rect 4844 11228 5124 11284
rect 4060 9774 4062 9826
rect 4114 9774 4116 9826
rect 4060 9762 4116 9774
rect 2940 8082 2996 8092
rect 3276 8036 3332 9212
rect 3500 9714 3668 9716
rect 3500 9662 3614 9714
rect 3666 9662 3668 9714
rect 3500 9660 3668 9662
rect 3500 8148 3556 9660
rect 3612 9650 3668 9660
rect 3948 9602 4004 9614
rect 3948 9550 3950 9602
rect 4002 9550 4004 9602
rect 3948 9154 4004 9550
rect 4172 9602 4228 9614
rect 4172 9550 4174 9602
rect 4226 9550 4228 9602
rect 4172 9492 4228 9550
rect 4172 9426 4228 9436
rect 3948 9102 3950 9154
rect 4002 9102 4004 9154
rect 3948 9090 4004 9102
rect 4284 9044 4340 10556
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4732 9940 4788 9950
rect 4732 9380 4788 9884
rect 4844 9938 4900 11228
rect 5180 11172 5236 11182
rect 5180 10722 5236 11116
rect 5180 10670 5182 10722
rect 5234 10670 5236 10722
rect 5180 10658 5236 10670
rect 5404 10610 5460 10622
rect 5404 10558 5406 10610
rect 5458 10558 5460 10610
rect 5292 10388 5348 10398
rect 5292 10294 5348 10332
rect 4956 10052 5012 10062
rect 5404 10052 5460 10558
rect 4956 9958 5012 9996
rect 5180 9996 5460 10052
rect 4844 9886 4846 9938
rect 4898 9886 4900 9938
rect 4844 9874 4900 9886
rect 4732 9314 4788 9324
rect 3948 8820 4004 8830
rect 3948 8258 4004 8764
rect 3948 8206 3950 8258
rect 4002 8206 4004 8258
rect 3948 8194 4004 8206
rect 3500 8082 3556 8092
rect 2828 7746 2884 7756
rect 3052 7980 3332 8036
rect 3724 8036 3780 8046
rect 2828 6580 2884 6590
rect 2884 6524 2996 6580
rect 2828 6486 2884 6524
rect 2716 6468 2772 6478
rect 2604 5794 2660 5806
rect 2604 5742 2606 5794
rect 2658 5742 2660 5794
rect 2604 5234 2660 5742
rect 2604 5182 2606 5234
rect 2658 5182 2660 5234
rect 2604 5170 2660 5182
rect 2268 5070 2270 5122
rect 2322 5070 2324 5122
rect 2268 5058 2324 5070
rect 2492 5012 2548 5022
rect 2492 4918 2548 4956
rect 2716 5010 2772 6412
rect 2716 4958 2718 5010
rect 2770 4958 2772 5010
rect 2716 4946 2772 4958
rect 2156 4498 2212 4508
rect 2828 4898 2884 4910
rect 2828 4846 2830 4898
rect 2882 4846 2884 4898
rect 2044 4286 2046 4338
rect 2098 4286 2100 4338
rect 2044 4274 2100 4286
rect 1036 3042 1092 3052
rect 2268 3442 2324 3454
rect 2268 3390 2270 3442
rect 2322 3390 2324 3442
rect 1148 2548 1204 2558
rect 1148 800 1204 2492
rect 2268 2548 2324 3390
rect 2828 3220 2884 4846
rect 2828 3154 2884 3164
rect 2940 2996 2996 6524
rect 3052 4226 3108 7980
rect 3724 7942 3780 7980
rect 3836 8034 3892 8046
rect 3836 7982 3838 8034
rect 3890 7982 3892 8034
rect 3500 7924 3556 7934
rect 3052 4174 3054 4226
rect 3106 4174 3108 4226
rect 3052 4162 3108 4174
rect 3276 6804 3332 6814
rect 3276 5012 3332 6748
rect 3500 5236 3556 7868
rect 3836 7588 3892 7982
rect 4060 8036 4116 8046
rect 4060 7942 4116 7980
rect 3948 7588 4004 7598
rect 3836 7586 4004 7588
rect 3836 7534 3950 7586
rect 4002 7534 4004 7586
rect 3836 7532 4004 7534
rect 3948 7522 4004 7532
rect 4172 7364 4228 7374
rect 4172 6802 4228 7308
rect 4172 6750 4174 6802
rect 4226 6750 4228 6802
rect 4172 6738 4228 6750
rect 3500 5170 3556 5180
rect 4172 6244 4228 6254
rect 3276 3780 3332 4956
rect 3276 3714 3332 3724
rect 3836 5010 3892 5022
rect 3836 4958 3838 5010
rect 3890 4958 3892 5010
rect 2268 2482 2324 2492
rect 2492 2940 2996 2996
rect 2492 800 2548 2940
rect 3836 2660 3892 4958
rect 4172 3666 4228 6188
rect 4284 5796 4340 8988
rect 4732 9044 4788 9054
rect 4732 9042 5012 9044
rect 4732 8990 4734 9042
rect 4786 8990 5012 9042
rect 4732 8988 5012 8990
rect 4732 8978 4788 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4732 8148 4788 8158
rect 4620 8146 4788 8148
rect 4620 8094 4734 8146
rect 4786 8094 4788 8146
rect 4620 8092 4788 8094
rect 4620 7252 4676 8092
rect 4732 8082 4788 8092
rect 4844 8034 4900 8046
rect 4844 7982 4846 8034
rect 4898 7982 4900 8034
rect 4844 7924 4900 7982
rect 4844 7858 4900 7868
rect 4732 7476 4788 7486
rect 4956 7476 5012 8988
rect 5180 8932 5236 9996
rect 5404 9716 5460 9726
rect 5404 9266 5460 9660
rect 5404 9214 5406 9266
rect 5458 9214 5460 9266
rect 5404 9202 5460 9214
rect 5180 8866 5236 8876
rect 5292 8930 5348 8942
rect 5292 8878 5294 8930
rect 5346 8878 5348 8930
rect 5292 8708 5348 8878
rect 5292 8642 5348 8652
rect 5068 8148 5124 8158
rect 5068 8054 5124 8092
rect 5516 7812 5572 11732
rect 5628 10948 5684 12238
rect 5740 11956 5796 11966
rect 5740 11862 5796 11900
rect 5852 11732 5908 14028
rect 5964 13188 6020 14254
rect 6076 14308 6132 14318
rect 6076 13412 6132 14252
rect 6412 14308 6468 15262
rect 6524 15316 6580 16046
rect 6524 15250 6580 15260
rect 6636 15148 6692 17836
rect 6748 17108 6804 20078
rect 6972 20188 7252 20244
rect 6748 17042 6804 17052
rect 6860 19572 6916 19582
rect 6972 19572 7028 20188
rect 7308 20132 7364 24558
rect 7420 23714 7476 23726
rect 7420 23662 7422 23714
rect 7474 23662 7476 23714
rect 7420 23492 7476 23662
rect 7532 23716 7588 25228
rect 7868 25282 7924 25294
rect 7868 25230 7870 25282
rect 7922 25230 7924 25282
rect 7644 24610 7700 24622
rect 7644 24558 7646 24610
rect 7698 24558 7700 24610
rect 7644 24500 7700 24558
rect 7644 24434 7700 24444
rect 7756 23716 7812 23726
rect 7532 23714 7812 23716
rect 7532 23662 7758 23714
rect 7810 23662 7812 23714
rect 7532 23660 7812 23662
rect 7420 23426 7476 23436
rect 7420 23156 7476 23166
rect 7420 23042 7476 23100
rect 7420 22990 7422 23042
rect 7474 22990 7476 23042
rect 7420 21924 7476 22990
rect 7420 21858 7476 21868
rect 7532 21476 7588 21486
rect 7532 21382 7588 21420
rect 7644 21028 7700 23660
rect 7756 23650 7812 23660
rect 7868 23604 7924 25230
rect 9548 25284 9604 25294
rect 8204 24612 8260 24622
rect 7868 23538 7924 23548
rect 8092 24610 8260 24612
rect 8092 24558 8206 24610
rect 8258 24558 8260 24610
rect 8092 24556 8260 24558
rect 8092 24498 8148 24556
rect 8204 24546 8260 24556
rect 8652 24612 8708 24622
rect 8652 24610 8820 24612
rect 8652 24558 8654 24610
rect 8706 24558 8820 24610
rect 8652 24556 8820 24558
rect 8652 24546 8708 24556
rect 8092 24446 8094 24498
rect 8146 24446 8148 24498
rect 7868 23044 7924 23054
rect 7868 22950 7924 22988
rect 8092 22932 8148 24446
rect 8764 24162 8820 24556
rect 9100 24610 9156 24622
rect 9100 24558 9102 24610
rect 9154 24558 9156 24610
rect 9100 24498 9156 24558
rect 9100 24446 9102 24498
rect 9154 24446 9156 24498
rect 9100 24434 9156 24446
rect 9548 24500 9604 25228
rect 9548 24434 9604 24444
rect 9996 24610 10052 24622
rect 9996 24558 9998 24610
rect 10050 24558 10052 24610
rect 9996 24276 10052 24558
rect 9996 24210 10052 24220
rect 10668 24610 10724 24622
rect 10668 24558 10670 24610
rect 10722 24558 10724 24610
rect 8764 24110 8766 24162
rect 8818 24110 8820 24162
rect 8764 24098 8820 24110
rect 9548 24162 9604 24174
rect 9548 24110 9550 24162
rect 9602 24110 9604 24162
rect 8652 24052 8708 24062
rect 8316 23828 8372 23838
rect 8316 23734 8372 23772
rect 8092 22866 8148 22876
rect 8204 23156 8260 23166
rect 7644 20962 7700 20972
rect 7756 22146 7812 22158
rect 7756 22094 7758 22146
rect 7810 22094 7812 22146
rect 7756 20692 7812 22094
rect 8092 22146 8148 22158
rect 8092 22094 8094 22146
rect 8146 22094 8148 22146
rect 7980 21812 8036 21822
rect 8092 21812 8148 22094
rect 7980 21810 8148 21812
rect 7980 21758 7982 21810
rect 8034 21758 8148 21810
rect 7980 21756 8148 21758
rect 7980 21746 8036 21756
rect 8092 21588 8148 21756
rect 8092 21522 8148 21532
rect 7756 20626 7812 20636
rect 7980 20692 8036 20702
rect 7980 20598 8036 20636
rect 7644 20580 7700 20590
rect 7644 20486 7700 20524
rect 7084 20076 7364 20132
rect 7868 20132 7924 20142
rect 8204 20132 8260 23100
rect 8540 23042 8596 23054
rect 8540 22990 8542 23042
rect 8594 22990 8596 23042
rect 8540 22932 8596 22990
rect 8540 22866 8596 22876
rect 8540 22148 8596 22158
rect 8540 22054 8596 22092
rect 8540 21474 8596 21486
rect 8540 21422 8542 21474
rect 8594 21422 8596 21474
rect 8540 21362 8596 21422
rect 8540 21310 8542 21362
rect 8594 21310 8596 21362
rect 8540 21298 8596 21310
rect 7084 19796 7140 20076
rect 7196 19908 7252 19918
rect 7252 19852 7476 19908
rect 7196 19776 7252 19852
rect 7084 19730 7140 19740
rect 6972 19516 7252 19572
rect 6860 16100 6916 19516
rect 7084 19348 7140 19358
rect 6972 17220 7028 17230
rect 6972 17106 7028 17164
rect 6972 17054 6974 17106
rect 7026 17054 7028 17106
rect 6972 17042 7028 17054
rect 7084 16884 7140 19292
rect 7196 18562 7252 19516
rect 7308 19458 7364 19470
rect 7308 19406 7310 19458
rect 7362 19406 7364 19458
rect 7308 18674 7364 19406
rect 7308 18622 7310 18674
rect 7362 18622 7364 18674
rect 7308 18610 7364 18622
rect 7196 18510 7198 18562
rect 7250 18510 7252 18562
rect 7196 18004 7252 18510
rect 7196 17938 7252 17948
rect 7196 17668 7252 17678
rect 7196 17574 7252 17612
rect 7420 17444 7476 19852
rect 7644 19906 7700 19918
rect 7644 19854 7646 19906
rect 7698 19854 7700 19906
rect 7644 19794 7700 19854
rect 7644 19742 7646 19794
rect 7698 19742 7700 19794
rect 7644 19458 7700 19742
rect 7644 19406 7646 19458
rect 7698 19406 7700 19458
rect 7644 19394 7700 19406
rect 7644 19124 7700 19134
rect 7644 19030 7700 19068
rect 7532 18450 7588 18462
rect 7532 18398 7534 18450
rect 7586 18398 7588 18450
rect 7532 18340 7588 18398
rect 7532 18274 7588 18284
rect 7532 17668 7588 17678
rect 7532 17574 7588 17612
rect 7420 17350 7476 17388
rect 7644 16996 7700 17006
rect 6860 16034 6916 16044
rect 6972 16828 7140 16884
rect 7420 16994 7700 16996
rect 7420 16942 7646 16994
rect 7698 16942 7700 16994
rect 7420 16940 7700 16942
rect 6748 15988 6804 15998
rect 6748 15876 6804 15932
rect 6860 15876 6916 15886
rect 6748 15874 6916 15876
rect 6748 15822 6862 15874
rect 6914 15822 6916 15874
rect 6748 15820 6916 15822
rect 6860 15810 6916 15820
rect 6972 15148 7028 16828
rect 7308 16100 7364 16110
rect 7084 15876 7140 15886
rect 7084 15782 7140 15820
rect 7196 15874 7252 15886
rect 7196 15822 7198 15874
rect 7250 15822 7252 15874
rect 7084 15428 7140 15438
rect 7196 15428 7252 15822
rect 7308 15652 7364 16044
rect 7308 15538 7364 15596
rect 7308 15486 7310 15538
rect 7362 15486 7364 15538
rect 7308 15474 7364 15486
rect 7420 15540 7476 16940
rect 7644 16930 7700 16940
rect 7756 16882 7812 16894
rect 7756 16830 7758 16882
rect 7810 16830 7812 16882
rect 7644 16660 7700 16670
rect 7420 15474 7476 15484
rect 7532 16658 7700 16660
rect 7532 16606 7646 16658
rect 7698 16606 7700 16658
rect 7532 16604 7700 16606
rect 7532 15538 7588 16604
rect 7644 16594 7700 16604
rect 7756 16324 7812 16830
rect 7756 16258 7812 16268
rect 7756 16100 7812 16110
rect 7868 16100 7924 20076
rect 8092 20076 8260 20132
rect 8316 21252 8372 21262
rect 8092 19460 8148 20076
rect 8092 19394 8148 19404
rect 8204 19906 8260 19918
rect 8204 19854 8206 19906
rect 8258 19854 8260 19906
rect 8204 19348 8260 19854
rect 8316 19794 8372 21196
rect 8540 20580 8596 20590
rect 8540 20486 8596 20524
rect 8316 19742 8318 19794
rect 8370 19742 8372 19794
rect 8316 19730 8372 19742
rect 8540 20020 8596 20030
rect 8204 19282 8260 19292
rect 8316 19460 8372 19470
rect 8092 19124 8148 19134
rect 8092 19030 8148 19068
rect 8204 19010 8260 19022
rect 8204 18958 8206 19010
rect 8258 18958 8260 19010
rect 8092 18676 8148 18686
rect 8092 18618 8148 18620
rect 8092 18566 8094 18618
rect 8146 18566 8148 18618
rect 8092 18554 8148 18566
rect 7980 18450 8036 18462
rect 7980 18398 7982 18450
rect 8034 18398 8036 18450
rect 7980 18228 8036 18398
rect 7980 18162 8036 18172
rect 8092 18226 8148 18238
rect 8092 18174 8094 18226
rect 8146 18174 8148 18226
rect 8092 17444 8148 18174
rect 8204 17668 8260 18958
rect 8316 18676 8372 19404
rect 8316 18610 8372 18620
rect 8540 18564 8596 19964
rect 8540 18498 8596 18508
rect 8652 18450 8708 23996
rect 9100 24052 9156 24062
rect 9100 23958 9156 23996
rect 8764 23492 8820 23502
rect 8764 22148 8820 23436
rect 9100 23042 9156 23054
rect 9100 22990 9102 23042
rect 9154 22990 9156 23042
rect 8988 22148 9044 22158
rect 8820 22146 9044 22148
rect 8820 22094 8990 22146
rect 9042 22094 9044 22146
rect 8820 22092 9044 22094
rect 8764 19460 8820 22092
rect 8988 22082 9044 22092
rect 9100 21812 9156 22990
rect 9548 23044 9604 24110
rect 9660 23714 9716 23726
rect 10108 23716 10164 23726
rect 9660 23662 9662 23714
rect 9714 23662 9716 23714
rect 9660 23604 9716 23662
rect 9660 23538 9716 23548
rect 9996 23714 10164 23716
rect 9996 23662 10110 23714
rect 10162 23662 10164 23714
rect 9996 23660 10164 23662
rect 9660 23044 9716 23054
rect 9548 23042 9716 23044
rect 9548 22990 9662 23042
rect 9714 22990 9716 23042
rect 9548 22988 9716 22990
rect 9100 21746 9156 21756
rect 9212 22260 9268 22270
rect 9100 21474 9156 21486
rect 9100 21422 9102 21474
rect 9154 21422 9156 21474
rect 8876 21362 8932 21374
rect 8876 21310 8878 21362
rect 8930 21310 8932 21362
rect 8876 19796 8932 21310
rect 8988 20916 9044 20926
rect 8988 20822 9044 20860
rect 9100 20580 9156 21422
rect 9100 20514 9156 20524
rect 9212 20356 9268 22204
rect 9548 22146 9604 22158
rect 9548 22094 9550 22146
rect 9602 22094 9604 22146
rect 9548 21700 9604 22094
rect 9660 22148 9716 22988
rect 9996 22372 10052 23660
rect 10108 23650 10164 23660
rect 10668 23268 10724 24558
rect 11116 24612 11172 24622
rect 11116 24518 11172 24556
rect 11228 24388 11284 24398
rect 11228 24050 11284 24332
rect 11228 23998 11230 24050
rect 11282 23998 11284 24050
rect 11228 23986 11284 23998
rect 11564 24388 11620 24398
rect 11452 23940 11508 23950
rect 10892 23714 10948 23726
rect 10892 23662 10894 23714
rect 10946 23662 10948 23714
rect 10892 23604 10948 23662
rect 10892 23538 10948 23548
rect 10668 23202 10724 23212
rect 10220 23156 10276 23166
rect 10220 23062 10276 23100
rect 9996 22306 10052 22316
rect 10668 23042 10724 23054
rect 11340 23044 11396 23054
rect 10668 22990 10670 23042
rect 10722 22990 10724 23042
rect 10668 22932 10724 22990
rect 10108 22260 10164 22270
rect 10108 22166 10164 22204
rect 10444 22148 10500 22158
rect 9660 22092 10052 22148
rect 9548 21634 9604 21644
rect 9772 21924 9828 21934
rect 9660 21474 9716 21486
rect 9660 21422 9662 21474
rect 9714 21422 9716 21474
rect 9660 21362 9716 21422
rect 9660 21310 9662 21362
rect 9714 21310 9716 21362
rect 9660 21298 9716 21310
rect 9772 21140 9828 21868
rect 9548 21084 9828 21140
rect 8876 19730 8932 19740
rect 8988 20300 9268 20356
rect 9324 20580 9380 20590
rect 8988 19906 9044 20300
rect 8988 19854 8990 19906
rect 9042 19854 9044 19906
rect 8764 19394 8820 19404
rect 8988 19122 9044 19854
rect 9212 20020 9268 20030
rect 8988 19070 8990 19122
rect 9042 19070 9044 19122
rect 8876 19012 8932 19022
rect 8652 18398 8654 18450
rect 8706 18398 8708 18450
rect 8428 17892 8484 17902
rect 8428 17798 8484 17836
rect 8204 17602 8260 17612
rect 8540 17556 8596 17566
rect 8540 17462 8596 17500
rect 8428 17444 8484 17454
rect 8092 17442 8484 17444
rect 8092 17390 8430 17442
rect 8482 17390 8484 17442
rect 8092 17388 8484 17390
rect 8428 17378 8484 17388
rect 8428 17220 8484 17230
rect 8428 17106 8484 17164
rect 8428 17054 8430 17106
rect 8482 17054 8484 17106
rect 8428 17042 8484 17054
rect 8540 17108 8596 17118
rect 8316 16996 8372 17006
rect 8204 16884 8260 16894
rect 8204 16790 8260 16828
rect 7532 15486 7534 15538
rect 7586 15486 7588 15538
rect 7532 15474 7588 15486
rect 7644 16098 7924 16100
rect 7644 16046 7758 16098
rect 7810 16046 7924 16098
rect 7644 16044 7924 16046
rect 8092 16660 8148 16670
rect 7084 15426 7252 15428
rect 7084 15374 7086 15426
rect 7138 15374 7252 15426
rect 7084 15372 7252 15374
rect 7084 15362 7140 15372
rect 6412 14242 6468 14252
rect 6524 15092 6692 15148
rect 6860 15092 7028 15148
rect 7084 15204 7140 15214
rect 6412 13860 6468 13870
rect 6524 13860 6580 15092
rect 6748 14306 6804 14318
rect 6748 14254 6750 14306
rect 6802 14254 6804 14306
rect 6412 13858 6580 13860
rect 6412 13806 6414 13858
rect 6466 13806 6580 13858
rect 6412 13804 6580 13806
rect 6636 14196 6692 14206
rect 6412 13794 6468 13804
rect 6300 13746 6356 13758
rect 6300 13694 6302 13746
rect 6354 13694 6356 13746
rect 6076 13356 6244 13412
rect 6076 13188 6132 13198
rect 5964 13186 6132 13188
rect 5964 13134 6078 13186
rect 6130 13134 6132 13186
rect 5964 13132 6132 13134
rect 6076 13122 6132 13132
rect 5964 12964 6020 12974
rect 6188 12964 6244 13356
rect 5964 12870 6020 12908
rect 6076 12908 6244 12964
rect 5740 11396 5796 11406
rect 5740 11302 5796 11340
rect 5628 10892 5796 10948
rect 5628 10724 5684 10734
rect 5628 10630 5684 10668
rect 5740 10612 5796 10892
rect 5740 10546 5796 10556
rect 5740 9714 5796 9726
rect 5740 9662 5742 9714
rect 5794 9662 5796 9714
rect 5740 9604 5796 9662
rect 5852 9716 5908 11676
rect 6076 11394 6132 12908
rect 6300 12292 6356 13694
rect 6412 13524 6468 13534
rect 6412 13430 6468 13468
rect 6636 13076 6692 14140
rect 6748 14084 6804 14254
rect 6748 14018 6804 14028
rect 6860 13412 6916 15092
rect 7084 14532 7140 15148
rect 7532 15204 7588 15242
rect 7532 15138 7588 15148
rect 7644 15092 7700 16044
rect 7756 16034 7812 16044
rect 7644 15026 7700 15036
rect 7756 15876 7812 15886
rect 6972 14476 7140 14532
rect 6972 13860 7028 14476
rect 7196 14418 7252 14430
rect 7196 14366 7198 14418
rect 7250 14366 7252 14418
rect 7196 14308 7252 14366
rect 7420 14420 7476 14430
rect 7196 14242 7252 14252
rect 7308 14306 7364 14318
rect 7308 14254 7310 14306
rect 7362 14254 7364 14306
rect 7308 14084 7364 14254
rect 7196 14028 7364 14084
rect 7084 13860 7140 13870
rect 6972 13858 7140 13860
rect 6972 13806 7086 13858
rect 7138 13806 7140 13858
rect 6972 13804 7140 13806
rect 7084 13794 7140 13804
rect 6412 13020 6692 13076
rect 6748 13356 6916 13412
rect 6412 12628 6468 13020
rect 6748 12964 6804 13356
rect 6412 12562 6468 12572
rect 6636 12908 6804 12964
rect 6860 13188 6916 13198
rect 6188 12236 6356 12292
rect 6188 11620 6244 12236
rect 6300 12068 6356 12078
rect 6300 11974 6356 12012
rect 6636 11620 6692 12908
rect 6748 12740 6804 12750
rect 6748 12402 6804 12684
rect 6748 12350 6750 12402
rect 6802 12350 6804 12402
rect 6748 11844 6804 12350
rect 6860 12404 6916 13132
rect 7196 13076 7252 14028
rect 7308 13860 7364 13870
rect 7308 13766 7364 13804
rect 7084 13020 7196 13076
rect 6972 12852 7028 12862
rect 6972 12758 7028 12796
rect 6972 12404 7028 12414
rect 6860 12402 7028 12404
rect 6860 12350 6974 12402
rect 7026 12350 7028 12402
rect 6860 12348 7028 12350
rect 6748 11778 6804 11788
rect 6860 12066 6916 12078
rect 6860 12014 6862 12066
rect 6914 12014 6916 12066
rect 6636 11564 6804 11620
rect 6188 11554 6244 11564
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 6076 11330 6132 11342
rect 6188 11396 6244 11406
rect 6412 11396 6468 11406
rect 6636 11396 6692 11406
rect 6188 11394 6356 11396
rect 6188 11342 6190 11394
rect 6242 11342 6356 11394
rect 6188 11340 6356 11342
rect 6188 11330 6244 11340
rect 6076 11170 6132 11182
rect 6076 11118 6078 11170
rect 6130 11118 6132 11170
rect 6076 10836 6132 11118
rect 6076 10770 6132 10780
rect 6188 10612 6244 10622
rect 6188 10518 6244 10556
rect 6188 10388 6244 10398
rect 6300 10388 6356 11340
rect 6412 11394 6580 11396
rect 6412 11342 6414 11394
rect 6466 11342 6580 11394
rect 6412 11340 6580 11342
rect 6412 11330 6468 11340
rect 6524 10836 6580 11340
rect 6636 11302 6692 11340
rect 6244 10332 6356 10388
rect 6412 10610 6468 10622
rect 6412 10558 6414 10610
rect 6466 10558 6468 10610
rect 6188 9826 6244 10332
rect 6412 10164 6468 10558
rect 6188 9774 6190 9826
rect 6242 9774 6244 9826
rect 5964 9716 6020 9726
rect 5852 9714 6020 9716
rect 5852 9662 5966 9714
rect 6018 9662 6020 9714
rect 5852 9660 6020 9662
rect 5964 9650 6020 9660
rect 5740 9538 5796 9548
rect 5852 9044 5908 9054
rect 5852 8950 5908 8988
rect 5964 8596 6020 8606
rect 5964 8370 6020 8540
rect 5964 8318 5966 8370
rect 6018 8318 6020 8370
rect 5964 8306 6020 8318
rect 6188 8258 6244 9774
rect 6300 10108 6468 10164
rect 6300 9716 6356 10108
rect 6412 9940 6468 9950
rect 6524 9940 6580 10780
rect 6636 11060 6692 11070
rect 6636 10834 6692 11004
rect 6636 10782 6638 10834
rect 6690 10782 6692 10834
rect 6636 10770 6692 10782
rect 6748 10724 6804 11564
rect 6860 10948 6916 12014
rect 6972 11844 7028 12348
rect 7084 12068 7140 13020
rect 7196 13010 7252 13020
rect 7308 13636 7364 13646
rect 7308 13074 7364 13580
rect 7420 13634 7476 14364
rect 7532 14306 7588 14318
rect 7532 14254 7534 14306
rect 7586 14254 7588 14306
rect 7532 14196 7588 14254
rect 7756 14196 7812 15820
rect 8092 15426 8148 16604
rect 8316 15538 8372 16940
rect 8540 16994 8596 17052
rect 8540 16942 8542 16994
rect 8594 16942 8596 16994
rect 8540 16930 8596 16942
rect 8652 16772 8708 18398
rect 8764 19010 8932 19012
rect 8764 18958 8878 19010
rect 8930 18958 8932 19010
rect 8764 18956 8932 18958
rect 8764 16996 8820 18956
rect 8876 18946 8932 18956
rect 8988 19012 9044 19070
rect 8988 18946 9044 18956
rect 9100 19348 9156 19358
rect 8876 18676 8932 18686
rect 9100 18676 9156 19292
rect 8876 18674 9156 18676
rect 8876 18622 8878 18674
rect 8930 18622 9156 18674
rect 8876 18620 9156 18622
rect 8876 18610 8932 18620
rect 9212 18564 9268 19964
rect 8988 18508 9268 18564
rect 8988 18450 9044 18508
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 18386 9044 18398
rect 9100 17778 9156 17790
rect 9100 17726 9102 17778
rect 9154 17726 9156 17778
rect 9100 17668 9156 17726
rect 9324 17668 9380 20524
rect 9436 20578 9492 20590
rect 9436 20526 9438 20578
rect 9490 20526 9492 20578
rect 9436 20020 9492 20526
rect 9436 19954 9492 19964
rect 9100 17612 9380 17668
rect 9212 17444 9268 17454
rect 9100 17108 9156 17118
rect 9100 17014 9156 17052
rect 8764 16930 8820 16940
rect 8652 16706 8708 16716
rect 8652 16436 8708 16446
rect 8316 15486 8318 15538
rect 8370 15486 8372 15538
rect 8316 15474 8372 15486
rect 8428 15986 8484 15998
rect 8428 15934 8430 15986
rect 8482 15934 8484 15986
rect 8428 15538 8484 15934
rect 8428 15486 8430 15538
rect 8482 15486 8484 15538
rect 8428 15474 8484 15486
rect 8092 15374 8094 15426
rect 8146 15374 8148 15426
rect 8092 15362 8148 15374
rect 8204 15316 8260 15326
rect 7980 14756 8036 14766
rect 7532 14140 7812 14196
rect 7420 13582 7422 13634
rect 7474 13582 7476 13634
rect 7420 13570 7476 13582
rect 7756 13524 7812 14140
rect 7868 14306 7924 14318
rect 7868 14254 7870 14306
rect 7922 14254 7924 14306
rect 7868 14084 7924 14254
rect 7868 14018 7924 14028
rect 7980 13972 8036 14700
rect 8204 14530 8260 15260
rect 8540 15314 8596 15326
rect 8540 15262 8542 15314
rect 8594 15262 8596 15314
rect 8540 15204 8596 15262
rect 8540 15138 8596 15148
rect 8204 14478 8206 14530
rect 8258 14478 8260 14530
rect 8204 14466 8260 14478
rect 8092 14308 8148 14318
rect 8092 14214 8148 14252
rect 8652 14308 8708 16380
rect 8988 16324 9044 16334
rect 8764 15540 8820 15550
rect 8764 15314 8820 15484
rect 8764 15262 8766 15314
rect 8818 15262 8820 15314
rect 8764 15250 8820 15262
rect 8988 15316 9044 16268
rect 8988 15250 9044 15260
rect 8764 14980 8820 14990
rect 8764 14642 8820 14924
rect 8764 14590 8766 14642
rect 8818 14590 8820 14642
rect 8764 14578 8820 14590
rect 8652 14242 8708 14252
rect 8092 13972 8148 13982
rect 7980 13970 8148 13972
rect 7980 13918 8094 13970
rect 8146 13918 8148 13970
rect 7980 13916 8148 13918
rect 8092 13906 8148 13916
rect 8876 13972 8932 13982
rect 8876 13878 8932 13916
rect 8204 13860 8260 13870
rect 8204 13766 8260 13804
rect 8764 13860 8820 13870
rect 8764 13766 8820 13804
rect 7868 13748 7924 13758
rect 7868 13654 7924 13692
rect 9100 13746 9156 13758
rect 9100 13694 9102 13746
rect 9154 13694 9156 13746
rect 7756 13468 8372 13524
rect 7308 13022 7310 13074
rect 7362 13022 7364 13074
rect 7308 13010 7364 13022
rect 8204 13076 8260 13086
rect 8204 12982 8260 13020
rect 7196 12738 7252 12750
rect 7196 12686 7198 12738
rect 7250 12686 7252 12738
rect 7196 12516 7252 12686
rect 7420 12740 7476 12750
rect 7420 12646 7476 12684
rect 7532 12738 7588 12750
rect 7532 12686 7534 12738
rect 7586 12686 7588 12738
rect 7532 12628 7588 12686
rect 7532 12562 7588 12572
rect 8092 12740 8148 12750
rect 7196 12450 7252 12460
rect 7532 12404 7588 12414
rect 7420 12178 7476 12190
rect 7420 12126 7422 12178
rect 7474 12126 7476 12178
rect 7084 12012 7364 12068
rect 6972 11778 7028 11788
rect 7196 11732 7252 11742
rect 6860 10882 6916 10892
rect 7084 11394 7140 11406
rect 7084 11342 7086 11394
rect 7138 11342 7140 11394
rect 6748 10668 6916 10724
rect 6748 10500 6804 10510
rect 6748 10406 6804 10444
rect 6412 9938 6580 9940
rect 6412 9886 6414 9938
rect 6466 9886 6580 9938
rect 6412 9884 6580 9886
rect 6412 9874 6468 9884
rect 6300 9660 6468 9716
rect 6412 9604 6468 9660
rect 6636 9714 6692 9726
rect 6636 9662 6638 9714
rect 6690 9662 6692 9714
rect 6412 9538 6468 9548
rect 6524 9602 6580 9614
rect 6524 9550 6526 9602
rect 6578 9550 6580 9602
rect 6524 9492 6580 9550
rect 6524 9426 6580 9436
rect 6524 9268 6580 9278
rect 6524 9174 6580 9212
rect 6412 9156 6468 9166
rect 6412 9062 6468 9100
rect 6300 9044 6356 9054
rect 6300 8950 6356 8988
rect 6636 8372 6692 9662
rect 6412 8316 6692 8372
rect 6860 8484 6916 10668
rect 7084 10052 7140 11342
rect 7196 10722 7252 11676
rect 7308 11506 7364 12012
rect 7308 11454 7310 11506
rect 7362 11454 7364 11506
rect 7308 11442 7364 11454
rect 7420 10834 7476 12126
rect 7532 11394 7588 12348
rect 7756 12292 7812 12302
rect 7532 11342 7534 11394
rect 7586 11342 7588 11394
rect 7532 11172 7588 11342
rect 7532 11106 7588 11116
rect 7644 11844 7700 11854
rect 7420 10782 7422 10834
rect 7474 10782 7476 10834
rect 7420 10770 7476 10782
rect 7196 10670 7198 10722
rect 7250 10670 7252 10722
rect 7196 10658 7252 10670
rect 7308 10724 7364 10734
rect 7084 9986 7140 9996
rect 7308 10050 7364 10668
rect 7532 10724 7588 10734
rect 7644 10724 7700 11788
rect 7756 11282 7812 12236
rect 7756 11230 7758 11282
rect 7810 11230 7812 11282
rect 7756 11172 7812 11230
rect 7980 12178 8036 12190
rect 7980 12126 7982 12178
rect 8034 12126 8036 12178
rect 7980 11284 8036 12126
rect 8092 12066 8148 12684
rect 8204 12404 8260 12414
rect 8316 12404 8372 13468
rect 9100 13188 9156 13694
rect 9100 13122 9156 13132
rect 8428 12964 8484 12974
rect 8428 12870 8484 12908
rect 8876 12852 8932 12862
rect 8764 12740 8820 12750
rect 8204 12402 8372 12404
rect 8204 12350 8206 12402
rect 8258 12350 8372 12402
rect 8204 12348 8372 12350
rect 8428 12738 8820 12740
rect 8428 12686 8766 12738
rect 8818 12686 8820 12738
rect 8428 12684 8820 12686
rect 8428 12402 8484 12684
rect 8764 12674 8820 12684
rect 8876 12516 8932 12796
rect 8428 12350 8430 12402
rect 8482 12350 8484 12402
rect 8204 12338 8260 12348
rect 8428 12338 8484 12350
rect 8540 12460 8932 12516
rect 8988 12628 9044 12638
rect 8092 12014 8094 12066
rect 8146 12014 8148 12066
rect 8092 12002 8148 12014
rect 8316 11732 8372 11742
rect 7980 11228 8260 11284
rect 7756 11116 8036 11172
rect 7532 10722 7700 10724
rect 7532 10670 7534 10722
rect 7586 10670 7700 10722
rect 7532 10668 7700 10670
rect 7532 10658 7588 10668
rect 7308 9998 7310 10050
rect 7362 9998 7364 10050
rect 7308 9986 7364 9998
rect 7420 10612 7476 10622
rect 7196 9380 7252 9390
rect 7084 9268 7140 9278
rect 7084 9174 7140 9212
rect 7196 9266 7252 9324
rect 7196 9214 7198 9266
rect 7250 9214 7252 9266
rect 7196 9202 7252 9214
rect 7308 9044 7364 9054
rect 7420 9044 7476 10556
rect 7756 10610 7812 10622
rect 7756 10558 7758 10610
rect 7810 10558 7812 10610
rect 7532 10500 7588 10510
rect 7532 9380 7588 10444
rect 7756 10052 7812 10558
rect 7756 9986 7812 9996
rect 7644 9828 7700 9838
rect 7644 9734 7700 9772
rect 7980 9828 8036 11116
rect 7980 9762 8036 9772
rect 8092 9940 8148 9950
rect 7868 9716 7924 9726
rect 7756 9714 7924 9716
rect 7756 9662 7870 9714
rect 7922 9662 7924 9714
rect 7756 9660 7924 9662
rect 7756 9380 7812 9660
rect 7868 9650 7924 9660
rect 7532 9324 7700 9380
rect 7532 9156 7588 9166
rect 7532 9062 7588 9100
rect 7308 9042 7476 9044
rect 7308 8990 7310 9042
rect 7362 8990 7476 9042
rect 7308 8988 7476 8990
rect 7308 8978 7364 8988
rect 6188 8206 6190 8258
rect 6242 8206 6244 8258
rect 5740 8146 5796 8158
rect 6188 8148 6244 8206
rect 6300 8260 6356 8270
rect 6300 8166 6356 8204
rect 5740 8094 5742 8146
rect 5794 8094 5796 8146
rect 5628 8036 5684 8046
rect 5628 7942 5684 7980
rect 5516 7756 5684 7812
rect 5516 7476 5572 7486
rect 4788 7420 5124 7476
rect 4732 7344 4788 7420
rect 4620 7196 5012 7252
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4620 6916 4676 6926
rect 4620 6356 4676 6860
rect 4732 6692 4788 6702
rect 4732 6598 4788 6636
rect 4844 6466 4900 6478
rect 4844 6414 4846 6466
rect 4898 6414 4900 6466
rect 4844 6356 4900 6414
rect 4620 6300 4900 6356
rect 4732 5796 4788 5806
rect 4284 5794 4788 5796
rect 4284 5742 4734 5794
rect 4786 5742 4788 5794
rect 4284 5740 4788 5742
rect 4732 5730 4788 5740
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4956 5460 5012 7196
rect 5068 6804 5124 7420
rect 5516 7382 5572 7420
rect 5068 6738 5124 6748
rect 5404 7250 5460 7262
rect 5404 7198 5406 7250
rect 5458 7198 5460 7250
rect 5068 6468 5124 6478
rect 5068 6466 5236 6468
rect 5068 6414 5070 6466
rect 5122 6414 5236 6466
rect 5068 6412 5236 6414
rect 5068 6402 5124 6412
rect 4476 5450 4740 5460
rect 4844 5404 5012 5460
rect 5068 6020 5124 6030
rect 4844 5236 4900 5404
rect 4732 5180 4900 5236
rect 4956 5236 5012 5246
rect 4732 4788 4788 5180
rect 4956 5142 5012 5180
rect 4732 4722 4788 4732
rect 4844 5012 4900 5022
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4172 3614 4174 3666
rect 4226 3614 4228 3666
rect 4172 3602 4228 3614
rect 4844 3666 4900 4956
rect 4956 4116 5012 4126
rect 4956 3778 5012 4060
rect 4956 3726 4958 3778
rect 5010 3726 5012 3778
rect 4956 3714 5012 3726
rect 4844 3614 4846 3666
rect 4898 3614 4900 3666
rect 4844 3602 4900 3614
rect 5068 3388 5124 5964
rect 5180 5908 5236 6412
rect 5180 5842 5236 5852
rect 5404 5460 5460 7198
rect 5628 6692 5684 7756
rect 5740 7476 5796 8094
rect 6076 8092 6244 8148
rect 5740 7420 6020 7476
rect 5964 7364 6020 7420
rect 5964 7298 6020 7308
rect 5628 6626 5684 6636
rect 5740 7250 5796 7262
rect 5740 7198 5742 7250
rect 5794 7198 5796 7250
rect 5740 6578 5796 7198
rect 6076 7252 6132 8092
rect 6412 7588 6468 8316
rect 6636 8146 6692 8158
rect 6636 8094 6638 8146
rect 6690 8094 6692 8146
rect 6636 8036 6692 8094
rect 6188 7532 6468 7588
rect 6524 7700 6580 7710
rect 6188 7474 6244 7532
rect 6188 7422 6190 7474
rect 6242 7422 6244 7474
rect 6188 7410 6244 7422
rect 6076 7196 6244 7252
rect 5964 7140 6020 7150
rect 5964 6802 6020 7084
rect 5964 6750 5966 6802
rect 6018 6750 6020 6802
rect 5964 6738 6020 6750
rect 6076 6804 6132 6814
rect 5740 6526 5742 6578
rect 5794 6526 5796 6578
rect 5628 6468 5684 6478
rect 5628 6374 5684 6412
rect 5516 6020 5572 6030
rect 5516 5926 5572 5964
rect 5404 5394 5460 5404
rect 5628 5236 5684 5246
rect 5740 5236 5796 6526
rect 5852 5348 5908 5358
rect 5852 5254 5908 5292
rect 5684 5180 5796 5236
rect 5628 5170 5684 5180
rect 5852 5124 5908 5134
rect 5740 5068 5852 5124
rect 5740 5010 5796 5068
rect 5852 5058 5908 5068
rect 5740 4958 5742 5010
rect 5794 4958 5796 5010
rect 5740 4946 5796 4958
rect 5964 4340 6020 4350
rect 6076 4340 6132 6748
rect 6188 6690 6244 7196
rect 6188 6638 6190 6690
rect 6242 6638 6244 6690
rect 6188 6020 6244 6638
rect 6188 5954 6244 5964
rect 6300 5236 6356 7532
rect 6412 7140 6468 7150
rect 6412 6690 6468 7084
rect 6412 6638 6414 6690
rect 6466 6638 6468 6690
rect 6412 6626 6468 6638
rect 6524 6692 6580 7644
rect 6636 7588 6692 7980
rect 6860 7700 6916 8428
rect 6860 7634 6916 7644
rect 7084 8932 7140 8942
rect 7084 8370 7140 8876
rect 7084 8318 7086 8370
rect 7138 8318 7140 8370
rect 7084 7698 7140 8318
rect 7084 7646 7086 7698
rect 7138 7646 7140 7698
rect 7084 7634 7140 7646
rect 7308 7700 7364 7710
rect 7308 7606 7364 7644
rect 6636 7522 6692 7532
rect 6860 7476 6916 7486
rect 6860 7382 6916 7420
rect 6972 7474 7028 7486
rect 6972 7422 6974 7474
rect 7026 7422 7028 7474
rect 6748 7364 6804 7374
rect 6636 6692 6692 6702
rect 6524 6690 6692 6692
rect 6524 6638 6638 6690
rect 6690 6638 6692 6690
rect 6524 6636 6692 6638
rect 6636 6626 6692 6636
rect 6748 5794 6804 7308
rect 6748 5742 6750 5794
rect 6802 5742 6804 5794
rect 6748 5730 6804 5742
rect 6860 6692 6916 6702
rect 6412 5236 6468 5246
rect 6300 5234 6468 5236
rect 6300 5182 6414 5234
rect 6466 5182 6468 5234
rect 6300 5180 6468 5182
rect 6412 5170 6468 5180
rect 6860 5124 6916 6636
rect 6972 5796 7028 7422
rect 7308 7476 7364 7486
rect 7308 6244 7364 7420
rect 7420 6802 7476 8988
rect 7644 8260 7700 9324
rect 7756 9314 7812 9324
rect 7868 9492 7924 9502
rect 7644 8204 7812 8260
rect 7644 8036 7700 8046
rect 7644 7942 7700 7980
rect 7420 6750 7422 6802
rect 7474 6750 7476 6802
rect 7420 6738 7476 6750
rect 7644 7252 7700 7262
rect 7532 6690 7588 6702
rect 7532 6638 7534 6690
rect 7586 6638 7588 6690
rect 7532 6580 7588 6638
rect 7532 6514 7588 6524
rect 7308 6178 7364 6188
rect 6972 5730 7028 5740
rect 7644 5794 7700 7196
rect 7644 5742 7646 5794
rect 7698 5742 7700 5794
rect 6636 4900 6692 4910
rect 5964 4338 6132 4340
rect 5964 4286 5966 4338
rect 6018 4286 6132 4338
rect 5964 4284 6132 4286
rect 6188 4676 6244 4686
rect 5964 4274 6020 4284
rect 5180 4228 5236 4238
rect 6188 4228 6244 4620
rect 6524 4452 6580 4462
rect 6524 4358 6580 4396
rect 5180 4226 5908 4228
rect 5180 4174 5182 4226
rect 5234 4174 5908 4226
rect 5180 4172 5908 4174
rect 5180 4162 5236 4172
rect 5852 3666 5908 4172
rect 5852 3614 5854 3666
rect 5906 3614 5908 3666
rect 5852 3602 5908 3614
rect 6076 4172 6244 4228
rect 5964 3556 6020 3566
rect 6076 3556 6132 4172
rect 5964 3554 6132 3556
rect 5964 3502 5966 3554
rect 6018 3502 6132 3554
rect 5964 3500 6132 3502
rect 6188 3780 6244 3790
rect 6188 3554 6244 3724
rect 6188 3502 6190 3554
rect 6242 3502 6244 3554
rect 5964 3490 6020 3500
rect 6188 3490 6244 3502
rect 6636 3388 6692 4844
rect 6748 4564 6804 4574
rect 6860 4564 6916 5068
rect 7644 5124 7700 5742
rect 7644 5058 7700 5068
rect 7420 5010 7476 5022
rect 7420 4958 7422 5010
rect 7474 4958 7476 5010
rect 7420 4900 7476 4958
rect 7420 4834 7476 4844
rect 6748 4562 6916 4564
rect 6748 4510 6750 4562
rect 6802 4510 6916 4562
rect 6748 4508 6916 4510
rect 6972 4564 7028 4574
rect 6748 4498 6804 4508
rect 6972 4470 7028 4508
rect 7644 4452 7700 4462
rect 7644 4358 7700 4396
rect 6860 4340 6916 4350
rect 6860 3778 6916 4284
rect 6860 3726 6862 3778
rect 6914 3726 6916 3778
rect 6860 3714 6916 3726
rect 7084 4114 7140 4126
rect 7084 4062 7086 4114
rect 7138 4062 7140 4114
rect 6748 3668 6804 3678
rect 6748 3574 6804 3612
rect 5068 3332 5236 3388
rect 3836 800 3892 2604
rect 5180 800 5236 3332
rect 6412 3332 6468 3342
rect 6412 3238 6468 3276
rect 6524 3332 6692 3388
rect 6524 800 6580 3332
rect 7084 2772 7140 4062
rect 7756 3388 7812 8204
rect 7868 6578 7924 9436
rect 7868 6526 7870 6578
rect 7922 6526 7924 6578
rect 7868 6514 7924 6526
rect 7980 7588 8036 7598
rect 7980 7140 8036 7532
rect 8092 7476 8148 9884
rect 8204 9604 8260 11228
rect 8316 11170 8372 11676
rect 8316 11118 8318 11170
rect 8370 11118 8372 11170
rect 8316 10388 8372 11118
rect 8428 10836 8484 10846
rect 8428 10742 8484 10780
rect 8316 10322 8372 10332
rect 8540 10164 8596 12460
rect 8540 10098 8596 10108
rect 8764 11956 8820 11966
rect 8428 9604 8484 9614
rect 8260 9602 8484 9604
rect 8260 9550 8430 9602
rect 8482 9550 8484 9602
rect 8260 9548 8484 9550
rect 8204 9472 8260 9548
rect 8428 9492 8484 9548
rect 8428 9426 8484 9436
rect 8316 9154 8372 9166
rect 8316 9102 8318 9154
rect 8370 9102 8372 9154
rect 8204 8820 8260 8830
rect 8204 8726 8260 8764
rect 8204 8484 8260 8494
rect 8204 8370 8260 8428
rect 8204 8318 8206 8370
rect 8258 8318 8260 8370
rect 8204 8306 8260 8318
rect 8316 8372 8372 9102
rect 8764 9154 8820 11900
rect 8988 11506 9044 12572
rect 9100 12404 9156 12414
rect 9100 12310 9156 12348
rect 8988 11454 8990 11506
rect 9042 11454 9044 11506
rect 8988 11442 9044 11454
rect 9212 11508 9268 17388
rect 9324 16324 9380 17612
rect 9436 19796 9492 19806
rect 9436 18452 9492 19740
rect 9436 16436 9492 18396
rect 9548 18340 9604 21084
rect 9884 20468 9940 20478
rect 9660 19906 9716 19918
rect 9660 19854 9662 19906
rect 9714 19854 9716 19906
rect 9660 19796 9716 19854
rect 9660 19236 9716 19740
rect 9884 19458 9940 20412
rect 9884 19406 9886 19458
rect 9938 19406 9940 19458
rect 9884 19394 9940 19406
rect 9772 19236 9828 19246
rect 9660 19234 9828 19236
rect 9660 19182 9774 19234
rect 9826 19182 9828 19234
rect 9660 19180 9828 19182
rect 9772 19170 9828 19180
rect 9884 19236 9940 19246
rect 9884 19122 9940 19180
rect 9884 19070 9886 19122
rect 9938 19070 9940 19122
rect 9884 19058 9940 19070
rect 9884 18676 9940 18686
rect 9884 18582 9940 18620
rect 9772 18564 9828 18574
rect 9772 18470 9828 18508
rect 9548 18284 9828 18340
rect 9660 18004 9716 18014
rect 9660 17444 9716 17948
rect 9660 17106 9716 17388
rect 9660 17054 9662 17106
rect 9714 17054 9716 17106
rect 9660 17042 9716 17054
rect 9436 16370 9492 16380
rect 9660 16660 9716 16670
rect 9324 16258 9380 16268
rect 9548 16212 9604 16222
rect 9324 15540 9380 15550
rect 9324 15148 9380 15484
rect 9548 15540 9604 16156
rect 9324 15092 9492 15148
rect 9324 14756 9380 14766
rect 9324 11844 9380 14700
rect 9324 11778 9380 11788
rect 9324 11620 9380 11630
rect 9324 11526 9380 11564
rect 9212 11442 9268 11452
rect 8876 11396 8932 11406
rect 8876 9940 8932 11340
rect 9100 11394 9156 11406
rect 9100 11342 9102 11394
rect 9154 11342 9156 11394
rect 9100 10836 9156 11342
rect 9100 10770 9156 10780
rect 9324 11060 9380 11070
rect 9436 11060 9492 15092
rect 9548 11394 9604 15484
rect 9660 14532 9716 16604
rect 9772 14756 9828 18284
rect 9884 18228 9940 18238
rect 9884 18134 9940 18172
rect 9772 14690 9828 14700
rect 9884 17556 9940 17566
rect 9996 17556 10052 22092
rect 10444 22054 10500 22092
rect 10668 22036 10724 22876
rect 11116 23042 11396 23044
rect 11116 22990 11342 23042
rect 11394 22990 11396 23042
rect 11116 22988 11396 22990
rect 11004 22148 11060 22158
rect 10668 21970 10724 21980
rect 10892 22146 11060 22148
rect 10892 22094 11006 22146
rect 11058 22094 11060 22146
rect 10892 22092 11060 22094
rect 10108 21812 10164 21822
rect 10108 21718 10164 21756
rect 10556 21812 10612 21822
rect 10556 21718 10612 21756
rect 10668 21700 10724 21710
rect 10220 20580 10276 20590
rect 10220 20486 10276 20524
rect 10668 20578 10724 21644
rect 10668 20526 10670 20578
rect 10722 20526 10724 20578
rect 10668 20244 10724 20526
rect 10444 20020 10500 20030
rect 10444 19926 10500 19964
rect 10444 19236 10500 19246
rect 10444 19142 10500 19180
rect 9940 17500 10052 17556
rect 10108 19124 10164 19134
rect 9660 14476 9828 14532
rect 9548 11342 9550 11394
rect 9602 11342 9604 11394
rect 9548 11330 9604 11342
rect 9660 14308 9716 14318
rect 9660 13074 9716 14252
rect 9772 13748 9828 14476
rect 9884 13972 9940 17500
rect 9996 15540 10052 15550
rect 9996 15426 10052 15484
rect 9996 15374 9998 15426
rect 10050 15374 10052 15426
rect 9996 15362 10052 15374
rect 10108 15426 10164 19068
rect 10668 19124 10724 20188
rect 10668 19058 10724 19068
rect 10780 21364 10836 21374
rect 10892 21364 10948 22092
rect 11004 22082 11060 22092
rect 11004 21924 11060 21934
rect 11004 21810 11060 21868
rect 11004 21758 11006 21810
rect 11058 21758 11060 21810
rect 11004 21746 11060 21758
rect 10780 21362 10948 21364
rect 10780 21310 10782 21362
rect 10834 21310 10948 21362
rect 10780 21308 10948 21310
rect 10780 18900 10836 21308
rect 10892 20132 10948 20142
rect 10892 20038 10948 20076
rect 10668 18844 10836 18900
rect 10892 19908 10948 19918
rect 10332 17668 10388 17678
rect 10332 17106 10388 17612
rect 10332 17054 10334 17106
rect 10386 17054 10388 17106
rect 10220 16996 10276 17006
rect 10220 16902 10276 16940
rect 10332 16772 10388 17054
rect 10556 16884 10612 16894
rect 10556 16790 10612 16828
rect 10108 15374 10110 15426
rect 10162 15374 10164 15426
rect 10108 15148 10164 15374
rect 9884 13906 9940 13916
rect 9996 15092 10164 15148
rect 10220 16716 10388 16772
rect 9996 14980 10052 15092
rect 9884 13748 9940 13758
rect 9772 13746 9940 13748
rect 9772 13694 9886 13746
rect 9938 13694 9940 13746
rect 9772 13692 9940 13694
rect 9884 13412 9940 13692
rect 9996 13636 10052 14924
rect 10220 14196 10276 16716
rect 10556 16210 10612 16222
rect 10556 16158 10558 16210
rect 10610 16158 10612 16210
rect 10332 15764 10388 15774
rect 10332 15538 10388 15708
rect 10332 15486 10334 15538
rect 10386 15486 10388 15538
rect 10332 15474 10388 15486
rect 10556 15540 10612 16158
rect 10556 15474 10612 15484
rect 10444 15316 10500 15326
rect 10108 14140 10276 14196
rect 10332 15204 10388 15214
rect 10108 13970 10164 14140
rect 10108 13918 10110 13970
rect 10162 13918 10164 13970
rect 10108 13860 10164 13918
rect 10220 13972 10276 13982
rect 10220 13878 10276 13916
rect 10332 13970 10388 15148
rect 10444 15148 10500 15260
rect 10444 15092 10612 15148
rect 10332 13918 10334 13970
rect 10386 13918 10388 13970
rect 10332 13906 10388 13918
rect 10108 13794 10164 13804
rect 10444 13746 10500 13758
rect 10444 13694 10446 13746
rect 10498 13694 10500 13746
rect 9996 13580 10164 13636
rect 9884 13346 9940 13356
rect 9660 13022 9662 13074
rect 9714 13022 9716 13074
rect 9660 11172 9716 13022
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 11844 9828 12126
rect 9772 11778 9828 11788
rect 9996 11844 10052 11854
rect 9884 11732 9940 11742
rect 9772 11508 9828 11518
rect 9772 11394 9828 11452
rect 9772 11342 9774 11394
rect 9826 11342 9828 11394
rect 9772 11330 9828 11342
rect 9772 11172 9828 11182
rect 9660 11116 9772 11172
rect 9772 11106 9828 11116
rect 9436 11004 9716 11060
rect 8988 10498 9044 10510
rect 8988 10446 8990 10498
rect 9042 10446 9044 10498
rect 8988 10164 9044 10446
rect 8988 10098 9044 10108
rect 8876 9884 9268 9940
rect 8988 9716 9044 9726
rect 8764 9102 8766 9154
rect 8818 9102 8820 9154
rect 8764 9090 8820 9102
rect 8876 9714 9044 9716
rect 8876 9662 8990 9714
rect 9042 9662 9044 9714
rect 8876 9660 9044 9662
rect 8540 9042 8596 9054
rect 8540 8990 8542 9042
rect 8594 8990 8596 9042
rect 8540 8932 8596 8990
rect 8540 8484 8596 8876
rect 8540 8418 8596 8428
rect 8876 8484 8932 9660
rect 8988 9650 9044 9660
rect 8876 8418 8932 8428
rect 8988 8820 9044 8830
rect 8316 8306 8372 8316
rect 8316 8036 8372 8046
rect 8204 7476 8260 7486
rect 8092 7474 8260 7476
rect 8092 7422 8206 7474
rect 8258 7422 8260 7474
rect 8092 7420 8260 7422
rect 8204 7410 8260 7420
rect 7980 5124 8036 7084
rect 8316 6580 8372 7980
rect 8764 8036 8820 8046
rect 8764 7942 8820 7980
rect 8876 8034 8932 8046
rect 8876 7982 8878 8034
rect 8930 7982 8932 8034
rect 8428 7812 8484 7822
rect 8428 7474 8484 7756
rect 8876 7700 8932 7982
rect 8876 7634 8932 7644
rect 8988 8034 9044 8764
rect 8988 7982 8990 8034
rect 9042 7982 9044 8034
rect 8428 7422 8430 7474
rect 8482 7422 8484 7474
rect 8428 7410 8484 7422
rect 8652 7252 8708 7262
rect 8652 7158 8708 7196
rect 8428 6580 8484 6590
rect 8316 6578 8484 6580
rect 8316 6526 8430 6578
rect 8482 6526 8484 6578
rect 8316 6524 8484 6526
rect 7868 5068 8036 5124
rect 8092 6244 8148 6254
rect 7868 3780 7924 5068
rect 7868 3714 7924 3724
rect 7196 3332 7812 3388
rect 7868 3444 7924 3482
rect 7868 3378 7924 3388
rect 7196 3220 7252 3332
rect 8092 3220 8148 6188
rect 8428 5234 8484 6524
rect 8876 6244 8932 6254
rect 8876 6018 8932 6188
rect 8876 5966 8878 6018
rect 8930 5966 8932 6018
rect 8876 5954 8932 5966
rect 8428 5182 8430 5234
rect 8482 5182 8484 5234
rect 8428 5012 8484 5182
rect 8428 4946 8484 4956
rect 8988 5012 9044 7982
rect 9100 7700 9156 7710
rect 9100 7606 9156 7644
rect 9212 6804 9268 9884
rect 9324 8258 9380 11004
rect 9660 10834 9716 11004
rect 9660 10782 9662 10834
rect 9714 10782 9716 10834
rect 9660 10770 9716 10782
rect 9772 10612 9828 10622
rect 9772 10518 9828 10556
rect 9772 9828 9828 9838
rect 9772 9734 9828 9772
rect 9548 9716 9604 9726
rect 9548 9622 9604 9660
rect 9884 9268 9940 11676
rect 9996 11172 10052 11788
rect 10108 11172 10164 13580
rect 10220 13412 10276 13422
rect 10220 12740 10276 13356
rect 10220 12066 10276 12684
rect 10220 12014 10222 12066
rect 10274 12014 10276 12066
rect 10220 11844 10276 12014
rect 10220 11778 10276 11788
rect 10220 11508 10276 11518
rect 10220 11396 10276 11452
rect 10220 11394 10388 11396
rect 10220 11342 10222 11394
rect 10274 11342 10388 11394
rect 10220 11340 10388 11342
rect 10220 11330 10276 11340
rect 10108 11116 10276 11172
rect 9996 11106 10052 11116
rect 9996 10836 10052 10846
rect 9996 10610 10052 10780
rect 9996 10558 9998 10610
rect 10050 10558 10052 10610
rect 9996 10546 10052 10558
rect 10220 10612 10276 11116
rect 10332 10836 10388 11340
rect 10444 11172 10500 13694
rect 10556 11394 10612 15092
rect 10668 11620 10724 18844
rect 10892 18676 10948 19852
rect 10892 18544 10948 18620
rect 11004 18564 11060 18574
rect 11004 18470 11060 18508
rect 10892 18228 10948 18238
rect 10892 18134 10948 18172
rect 11116 16996 11172 22988
rect 11340 22978 11396 22988
rect 11340 22484 11396 22494
rect 11452 22484 11508 23884
rect 11396 22428 11508 22484
rect 11340 22352 11396 22428
rect 11452 21474 11508 21486
rect 11452 21422 11454 21474
rect 11506 21422 11508 21474
rect 11452 21362 11508 21422
rect 11452 21310 11454 21362
rect 11506 21310 11508 21362
rect 11452 21298 11508 21310
rect 11564 20916 11620 24332
rect 12236 24052 12292 24062
rect 12236 23958 12292 23996
rect 13468 24052 13524 25340
rect 14476 24388 14532 24398
rect 13468 23986 13524 23996
rect 14028 24164 14084 24174
rect 14028 24050 14084 24108
rect 14028 23998 14030 24050
rect 14082 23998 14084 24050
rect 14028 23986 14084 23998
rect 14476 24050 14532 24332
rect 14476 23998 14478 24050
rect 14530 23998 14532 24050
rect 14476 23986 14532 23998
rect 15036 24052 15092 24062
rect 15036 23958 15092 23996
rect 13580 23940 13636 23950
rect 13580 23846 13636 23884
rect 11900 23714 11956 23726
rect 11900 23662 11902 23714
rect 11954 23662 11956 23714
rect 11452 20578 11508 20590
rect 11452 20526 11454 20578
rect 11506 20526 11508 20578
rect 11340 20244 11396 20254
rect 11340 20150 11396 20188
rect 11340 19458 11396 19470
rect 11340 19406 11342 19458
rect 11394 19406 11396 19458
rect 11228 19010 11284 19022
rect 11228 18958 11230 19010
rect 11282 18958 11284 19010
rect 11228 18676 11284 18958
rect 11228 18610 11284 18620
rect 11228 17556 11284 17566
rect 11228 17462 11284 17500
rect 11004 16940 11172 16996
rect 11340 16994 11396 19406
rect 11340 16942 11342 16994
rect 11394 16942 11396 16994
rect 10892 16772 10948 16782
rect 10892 15426 10948 16716
rect 10892 15374 10894 15426
rect 10946 15374 10948 15426
rect 10780 15314 10836 15326
rect 10780 15262 10782 15314
rect 10834 15262 10836 15314
rect 10780 14980 10836 15262
rect 10892 15316 10948 15374
rect 10892 15250 10948 15260
rect 10780 14914 10836 14924
rect 10892 14418 10948 14430
rect 10892 14366 10894 14418
rect 10946 14366 10948 14418
rect 10892 13972 10948 14366
rect 10892 13906 10948 13916
rect 11004 12516 11060 16940
rect 11228 16884 11284 16894
rect 11116 15986 11172 15998
rect 11116 15934 11118 15986
rect 11170 15934 11172 15986
rect 11116 15764 11172 15934
rect 11228 15986 11284 16828
rect 11340 16660 11396 16942
rect 11340 16594 11396 16604
rect 11452 18228 11508 20526
rect 11564 19458 11620 20860
rect 11564 19406 11566 19458
rect 11618 19406 11620 19458
rect 11564 19236 11620 19406
rect 11676 23604 11732 23614
rect 11676 19460 11732 23548
rect 11900 23604 11956 23662
rect 11900 23538 11956 23548
rect 12684 23716 12740 23726
rect 12012 23044 12068 23054
rect 12012 23042 12180 23044
rect 12012 22990 12014 23042
rect 12066 22990 12180 23042
rect 12012 22988 12180 22990
rect 12012 22978 12068 22988
rect 11788 22146 11844 22158
rect 11788 22094 11790 22146
rect 11842 22094 11844 22146
rect 11788 21812 11844 22094
rect 11788 21746 11844 21756
rect 12012 21476 12068 21486
rect 12012 21382 12068 21420
rect 11900 20916 11956 20926
rect 11900 20822 11956 20860
rect 12124 20804 12180 22988
rect 12460 23042 12516 23054
rect 12460 22990 12462 23042
rect 12514 22990 12516 23042
rect 12124 20738 12180 20748
rect 12236 22820 12292 22830
rect 12012 19908 12068 19918
rect 11676 19394 11732 19404
rect 11900 19852 12012 19908
rect 11676 19236 11732 19246
rect 11564 19234 11732 19236
rect 11564 19182 11678 19234
rect 11730 19182 11732 19234
rect 11564 19180 11732 19182
rect 11676 19170 11732 19180
rect 11788 18788 11844 18798
rect 11788 18674 11844 18732
rect 11788 18622 11790 18674
rect 11842 18622 11844 18674
rect 11788 18610 11844 18622
rect 11900 18564 11956 19852
rect 12012 19776 12068 19852
rect 12236 19458 12292 22764
rect 12348 22148 12404 22158
rect 12348 22054 12404 22092
rect 12348 21924 12404 21934
rect 12348 21474 12404 21868
rect 12348 21422 12350 21474
rect 12402 21422 12404 21474
rect 12348 21362 12404 21422
rect 12348 21310 12350 21362
rect 12402 21310 12404 21362
rect 12348 21298 12404 21310
rect 12460 20804 12516 22990
rect 12684 23044 12740 23660
rect 13020 23156 13076 23166
rect 13020 23062 13076 23100
rect 14028 23156 14084 23166
rect 12684 22148 12740 22988
rect 13468 23042 13524 23054
rect 13468 22990 13470 23042
rect 13522 22990 13524 23042
rect 13468 22932 13524 22990
rect 13804 23044 13860 23054
rect 13804 22950 13860 22988
rect 13468 22866 13524 22876
rect 14028 22260 14084 23100
rect 12684 22082 12740 22092
rect 12908 22146 12964 22158
rect 12908 22094 12910 22146
rect 12962 22094 12964 22146
rect 12908 21924 12964 22094
rect 12908 21858 12964 21868
rect 13132 22148 13188 22158
rect 12348 20748 12516 20804
rect 12908 20804 12964 20814
rect 12348 20020 12404 20748
rect 12460 20580 12516 20590
rect 12460 20486 12516 20524
rect 12908 20578 12964 20748
rect 12908 20526 12910 20578
rect 12962 20526 12964 20578
rect 12908 20244 12964 20526
rect 12908 20178 12964 20188
rect 12460 20132 12516 20142
rect 12460 20038 12516 20076
rect 12348 19954 12404 19964
rect 13020 19906 13076 19918
rect 13020 19854 13022 19906
rect 13074 19854 13076 19906
rect 12236 19406 12238 19458
rect 12290 19406 12292 19458
rect 12236 19236 12292 19406
rect 12124 19180 12292 19236
rect 12572 19460 12628 19470
rect 11900 18498 11956 18508
rect 12012 19012 12068 19022
rect 11452 16212 11508 18172
rect 12012 17666 12068 18956
rect 12124 18674 12180 19180
rect 12236 19010 12292 19022
rect 12236 18958 12238 19010
rect 12290 18958 12292 19010
rect 12236 18788 12292 18958
rect 12236 18732 12516 18788
rect 12124 18622 12126 18674
rect 12178 18622 12180 18674
rect 12124 18610 12180 18622
rect 12236 18564 12292 18574
rect 12012 17614 12014 17666
rect 12066 17614 12068 17666
rect 11676 17556 11732 17566
rect 11564 17220 11620 17230
rect 11564 17106 11620 17164
rect 11564 17054 11566 17106
rect 11618 17054 11620 17106
rect 11564 17042 11620 17054
rect 11676 17106 11732 17500
rect 11676 17054 11678 17106
rect 11730 17054 11732 17106
rect 11676 17042 11732 17054
rect 11900 16996 11956 17006
rect 11900 16902 11956 16940
rect 11788 16884 11844 16894
rect 11788 16790 11844 16828
rect 12012 16660 12068 17614
rect 12124 17668 12180 17678
rect 12124 16772 12180 17612
rect 12124 16706 12180 16716
rect 11228 15934 11230 15986
rect 11282 15934 11284 15986
rect 11228 15922 11284 15934
rect 11340 16156 11508 16212
rect 11788 16604 12068 16660
rect 12236 16660 12292 18508
rect 11340 15764 11396 16156
rect 11452 15988 11508 15998
rect 11452 15894 11508 15932
rect 11116 15698 11172 15708
rect 11228 15708 11396 15764
rect 11116 15316 11172 15326
rect 11116 15222 11172 15260
rect 11228 14308 11284 15708
rect 11676 15426 11732 15438
rect 11676 15374 11678 15426
rect 11730 15374 11732 15426
rect 11564 15316 11620 15326
rect 11564 15222 11620 15260
rect 11676 14756 11732 15374
rect 11676 14690 11732 14700
rect 11788 15092 11844 16604
rect 12236 16594 12292 16604
rect 12348 18228 12404 18238
rect 12124 16212 12180 16222
rect 11900 15988 11956 15998
rect 11900 15894 11956 15932
rect 12012 15876 12068 15886
rect 12012 15782 12068 15820
rect 11900 15540 11956 15550
rect 11900 15446 11956 15484
rect 11228 14242 11284 14252
rect 11564 14532 11620 14542
rect 11788 14532 11844 15036
rect 12124 15428 12180 16156
rect 12124 14644 12180 15372
rect 12236 15874 12292 15886
rect 12236 15822 12238 15874
rect 12290 15822 12292 15874
rect 12236 15314 12292 15822
rect 12236 15262 12238 15314
rect 12290 15262 12292 15314
rect 12236 15250 12292 15262
rect 12236 14644 12292 14654
rect 12124 14642 12292 14644
rect 12124 14590 12238 14642
rect 12290 14590 12292 14642
rect 12124 14588 12292 14590
rect 12236 14578 12292 14588
rect 11564 14530 11844 14532
rect 11564 14478 11566 14530
rect 11618 14478 11844 14530
rect 11564 14476 11844 14478
rect 11116 14084 11172 14094
rect 11116 13970 11172 14028
rect 11116 13918 11118 13970
rect 11170 13918 11172 13970
rect 11116 13906 11172 13918
rect 11564 13524 11620 14476
rect 11788 14308 11844 14318
rect 11788 13970 11844 14252
rect 11788 13918 11790 13970
rect 11842 13918 11844 13970
rect 11788 13906 11844 13918
rect 12012 14084 12068 14094
rect 12012 13970 12068 14028
rect 12012 13918 12014 13970
rect 12066 13918 12068 13970
rect 12012 13906 12068 13918
rect 11564 13458 11620 13468
rect 11676 13748 11732 13758
rect 12348 13748 12404 18172
rect 12460 17668 12516 18732
rect 12460 17602 12516 17612
rect 12572 16994 12628 19404
rect 12796 19458 12852 19470
rect 12796 19406 12798 19458
rect 12850 19406 12852 19458
rect 12684 19012 12740 19022
rect 12684 18918 12740 18956
rect 12684 18788 12740 18798
rect 12684 18562 12740 18732
rect 12796 18676 12852 19406
rect 12796 18674 12964 18676
rect 12796 18622 12798 18674
rect 12850 18622 12964 18674
rect 12796 18620 12964 18622
rect 12796 18610 12852 18620
rect 12684 18510 12686 18562
rect 12738 18510 12740 18562
rect 12684 18498 12740 18510
rect 12908 18340 12964 18620
rect 12908 18274 12964 18284
rect 12796 18228 12852 18238
rect 12796 18134 12852 18172
rect 13020 18004 13076 19854
rect 13020 17938 13076 17948
rect 12684 17668 12740 17706
rect 12684 17602 12740 17612
rect 12908 17556 12964 17566
rect 12684 17442 12740 17454
rect 12684 17390 12686 17442
rect 12738 17390 12740 17442
rect 12684 17220 12740 17390
rect 12684 17154 12740 17164
rect 12796 17444 12852 17454
rect 12572 16942 12574 16994
rect 12626 16942 12628 16994
rect 12572 16930 12628 16942
rect 12684 16996 12740 17006
rect 12796 16996 12852 17388
rect 12684 16994 12852 16996
rect 12684 16942 12686 16994
rect 12738 16942 12852 16994
rect 12684 16940 12852 16942
rect 12684 16930 12740 16940
rect 12796 16772 12852 16940
rect 12796 16706 12852 16716
rect 12572 16660 12628 16670
rect 12572 15652 12628 16604
rect 12684 16658 12740 16670
rect 12684 16606 12686 16658
rect 12738 16606 12740 16658
rect 12684 16548 12740 16606
rect 12908 16548 12964 17500
rect 12740 16492 12964 16548
rect 12684 16482 12740 16492
rect 12796 16324 12852 16334
rect 12796 16230 12852 16268
rect 12684 15986 12740 15998
rect 12684 15934 12686 15986
rect 12738 15934 12740 15986
rect 12684 15764 12740 15934
rect 12684 15698 12740 15708
rect 12796 15988 12852 15998
rect 12572 15538 12628 15596
rect 12572 15486 12574 15538
rect 12626 15486 12628 15538
rect 12572 15474 12628 15486
rect 12796 15538 12852 15932
rect 12796 15486 12798 15538
rect 12850 15486 12852 15538
rect 12796 15474 12852 15486
rect 12908 15764 12964 15774
rect 12684 15316 12740 15326
rect 12460 15204 12516 15242
rect 12460 15138 12516 15148
rect 12684 14530 12740 15260
rect 12684 14478 12686 14530
rect 12738 14478 12740 14530
rect 12684 14466 12740 14478
rect 12572 14420 12628 14430
rect 12460 13972 12516 13982
rect 12460 13858 12516 13916
rect 12572 13970 12628 14364
rect 12796 14420 12852 14430
rect 12908 14420 12964 15708
rect 13020 15428 13076 15438
rect 13020 14530 13076 15372
rect 13020 14478 13022 14530
rect 13074 14478 13076 14530
rect 13020 14466 13076 14478
rect 12796 14418 12964 14420
rect 12796 14366 12798 14418
rect 12850 14366 12964 14418
rect 12796 14364 12964 14366
rect 12796 14354 12852 14364
rect 12572 13918 12574 13970
rect 12626 13918 12628 13970
rect 12572 13906 12628 13918
rect 12460 13806 12462 13858
rect 12514 13806 12516 13858
rect 12460 13794 12516 13806
rect 12796 13860 12852 13870
rect 12796 13766 12852 13804
rect 11676 13746 12404 13748
rect 11676 13694 11678 13746
rect 11730 13694 12404 13746
rect 11676 13692 12404 13694
rect 11004 12460 11172 12516
rect 11004 12292 11060 12302
rect 11004 12198 11060 12236
rect 10892 11956 10948 11966
rect 10892 11954 11060 11956
rect 10892 11902 10894 11954
rect 10946 11902 11060 11954
rect 10892 11900 11060 11902
rect 10892 11890 10948 11900
rect 10780 11620 10836 11630
rect 10724 11618 10836 11620
rect 10724 11566 10782 11618
rect 10834 11566 10836 11618
rect 10724 11564 10836 11566
rect 10668 11488 10724 11564
rect 10556 11342 10558 11394
rect 10610 11342 10612 11394
rect 10556 11330 10612 11342
rect 10668 11172 10724 11182
rect 10444 11170 10724 11172
rect 10444 11118 10670 11170
rect 10722 11118 10724 11170
rect 10444 11116 10724 11118
rect 10668 11106 10724 11116
rect 10332 10780 10724 10836
rect 10668 10722 10724 10780
rect 10668 10670 10670 10722
rect 10722 10670 10724 10722
rect 10668 10658 10724 10670
rect 10332 10612 10388 10622
rect 10220 10610 10388 10612
rect 10220 10558 10334 10610
rect 10386 10558 10388 10610
rect 10220 10556 10388 10558
rect 10332 10546 10388 10556
rect 10220 10388 10276 10426
rect 10220 10322 10276 10332
rect 10780 10388 10836 11564
rect 11004 11394 11060 11900
rect 11004 11342 11006 11394
rect 11058 11342 11060 11394
rect 11004 10836 11060 11342
rect 11004 10770 11060 10780
rect 10780 10322 10836 10332
rect 10220 10164 10276 10174
rect 10108 10050 10164 10062
rect 10108 9998 10110 10050
rect 10162 9998 10164 10050
rect 9996 9604 10052 9614
rect 9996 9510 10052 9548
rect 9996 9268 10052 9278
rect 9884 9266 10052 9268
rect 9884 9214 9998 9266
rect 10050 9214 10052 9266
rect 9884 9212 10052 9214
rect 9996 9202 10052 9212
rect 10108 9266 10164 9998
rect 10220 9826 10276 10108
rect 11116 9828 11172 12460
rect 11564 12292 11620 12302
rect 11228 11396 11284 11406
rect 11228 11302 11284 11340
rect 11452 11396 11508 11406
rect 11228 10612 11284 10622
rect 11228 10518 11284 10556
rect 11340 10388 11396 10398
rect 11340 10294 11396 10332
rect 10220 9774 10222 9826
rect 10274 9774 10276 9826
rect 10220 9762 10276 9774
rect 11004 9772 11172 9828
rect 10108 9214 10110 9266
rect 10162 9214 10164 9266
rect 10108 9202 10164 9214
rect 10780 9716 10836 9726
rect 9884 9042 9940 9054
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9324 8206 9326 8258
rect 9378 8206 9380 8258
rect 9324 7252 9380 8206
rect 9324 7186 9380 7196
rect 9548 8820 9604 8830
rect 8988 4676 9044 4956
rect 8988 4610 9044 4620
rect 9100 6748 9268 6804
rect 9324 7028 9380 7038
rect 8988 4228 9044 4238
rect 9100 4228 9156 6748
rect 9212 6578 9268 6590
rect 9212 6526 9214 6578
rect 9266 6526 9268 6578
rect 9212 5684 9268 6526
rect 9324 6578 9380 6972
rect 9548 6690 9604 8764
rect 9884 7700 9940 8990
rect 10108 9044 10164 9054
rect 9996 8260 10052 8270
rect 9996 8166 10052 8204
rect 9884 7634 9940 7644
rect 9772 7362 9828 7374
rect 9772 7310 9774 7362
rect 9826 7310 9828 7362
rect 9772 6916 9828 7310
rect 9772 6850 9828 6860
rect 9996 7252 10052 7262
rect 9548 6638 9550 6690
rect 9602 6638 9604 6690
rect 9548 6626 9604 6638
rect 9996 6690 10052 7196
rect 9996 6638 9998 6690
rect 10050 6638 10052 6690
rect 9996 6626 10052 6638
rect 9324 6526 9326 6578
rect 9378 6526 9380 6578
rect 9324 6514 9380 6526
rect 9996 6468 10052 6478
rect 9884 6132 9940 6142
rect 9884 5906 9940 6076
rect 9884 5854 9886 5906
rect 9938 5854 9940 5906
rect 9884 5842 9940 5854
rect 9996 5906 10052 6412
rect 10108 6132 10164 8988
rect 10444 9042 10500 9054
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 8932 10500 8990
rect 10444 8596 10500 8876
rect 10780 8820 10836 9660
rect 10780 8754 10836 8764
rect 10892 9604 10948 9614
rect 10892 8708 10948 9548
rect 10892 8642 10948 8652
rect 11004 9156 11060 9772
rect 11116 9604 11172 9614
rect 11116 9602 11284 9604
rect 11116 9550 11118 9602
rect 11170 9550 11284 9602
rect 11116 9548 11284 9550
rect 11116 9538 11172 9548
rect 11116 9156 11172 9166
rect 11004 9154 11172 9156
rect 11004 9102 11118 9154
rect 11170 9102 11172 9154
rect 11004 9100 11172 9102
rect 10444 8530 10500 8540
rect 10332 8484 10388 8494
rect 10332 6690 10388 8428
rect 10668 8146 10724 8158
rect 10668 8094 10670 8146
rect 10722 8094 10724 8146
rect 10332 6638 10334 6690
rect 10386 6638 10388 6690
rect 10332 6626 10388 6638
rect 10444 7586 10500 7598
rect 10444 7534 10446 7586
rect 10498 7534 10500 7586
rect 10444 6690 10500 7534
rect 10556 7476 10612 7486
rect 10556 7382 10612 7420
rect 10668 7362 10724 8094
rect 10780 7700 10836 7710
rect 10780 7606 10836 7644
rect 11004 7698 11060 9100
rect 11116 9090 11172 9100
rect 11228 8708 11284 9548
rect 11228 8642 11284 8652
rect 11004 7646 11006 7698
rect 11058 7646 11060 7698
rect 10668 7310 10670 7362
rect 10722 7310 10724 7362
rect 10668 7298 10724 7310
rect 11004 7252 11060 7646
rect 11004 7186 11060 7196
rect 11228 8260 11284 8270
rect 10444 6638 10446 6690
rect 10498 6638 10500 6690
rect 10444 6626 10500 6638
rect 10556 7140 10612 7150
rect 10556 6690 10612 7084
rect 10556 6638 10558 6690
rect 10610 6638 10612 6690
rect 10556 6626 10612 6638
rect 11228 6804 11284 8204
rect 11116 6468 11172 6478
rect 11004 6466 11172 6468
rect 11004 6414 11118 6466
rect 11170 6414 11172 6466
rect 11004 6412 11172 6414
rect 10332 6132 10388 6142
rect 10108 6130 10388 6132
rect 10108 6078 10334 6130
rect 10386 6078 10388 6130
rect 10108 6076 10388 6078
rect 10332 6066 10388 6076
rect 9996 5854 9998 5906
rect 10050 5854 10052 5906
rect 9212 5618 9268 5628
rect 9884 4788 9940 4798
rect 9772 4676 9828 4686
rect 9772 4562 9828 4620
rect 9772 4510 9774 4562
rect 9826 4510 9828 4562
rect 9772 4498 9828 4510
rect 8988 4226 9100 4228
rect 8988 4174 8990 4226
rect 9042 4174 9100 4226
rect 8988 4172 9100 4174
rect 8988 4162 9044 4172
rect 9100 4096 9156 4172
rect 9212 4452 9268 4462
rect 8876 3780 8932 3790
rect 8876 3666 8932 3724
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 8876 3602 8932 3614
rect 7196 3154 7252 3164
rect 7868 3164 8148 3220
rect 7084 2706 7140 2716
rect 7868 800 7924 3164
rect 9212 800 9268 4396
rect 9884 4450 9940 4732
rect 9884 4398 9886 4450
rect 9938 4398 9940 4450
rect 9884 4386 9940 4398
rect 9996 4116 10052 5854
rect 10220 5906 10276 5918
rect 10220 5854 10222 5906
rect 10274 5854 10276 5906
rect 10108 5794 10164 5806
rect 10108 5742 10110 5794
rect 10162 5742 10164 5794
rect 10108 5348 10164 5742
rect 10220 5796 10276 5854
rect 10220 5730 10276 5740
rect 11004 5906 11060 6412
rect 11116 6402 11172 6412
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5348 11060 5854
rect 10108 5292 10612 5348
rect 10556 5234 10612 5292
rect 11004 5282 11060 5292
rect 10556 5182 10558 5234
rect 10610 5182 10612 5234
rect 10556 5170 10612 5182
rect 9996 4050 10052 4060
rect 10108 5124 10164 5134
rect 10108 3778 10164 5068
rect 11228 5122 11284 6748
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 10556 4452 10612 4462
rect 10556 4338 10612 4396
rect 11228 4452 11284 5070
rect 11228 4386 11284 4396
rect 11452 5796 11508 11340
rect 11564 10948 11620 12236
rect 11676 12068 11732 13692
rect 12460 13524 12516 13534
rect 12460 12964 12516 13468
rect 12684 13524 12740 13534
rect 12572 12964 12628 12974
rect 12460 12962 12628 12964
rect 12460 12910 12574 12962
rect 12626 12910 12628 12962
rect 12460 12908 12628 12910
rect 11788 12852 11844 12862
rect 11788 12850 12516 12852
rect 11788 12798 11790 12850
rect 11842 12798 12516 12850
rect 11788 12796 12516 12798
rect 11788 12786 11844 12796
rect 11676 12002 11732 12012
rect 12236 11844 12292 11854
rect 12236 11394 12292 11788
rect 12460 11508 12516 12796
rect 12572 12068 12628 12908
rect 12572 12002 12628 12012
rect 12572 11508 12628 11518
rect 12460 11506 12628 11508
rect 12460 11454 12574 11506
rect 12626 11454 12628 11506
rect 12460 11452 12628 11454
rect 12572 11442 12628 11452
rect 12236 11342 12238 11394
rect 12290 11342 12292 11394
rect 12236 11330 12292 11342
rect 12684 11394 12740 13468
rect 12684 11342 12686 11394
rect 12738 11342 12740 11394
rect 12684 11330 12740 11342
rect 12908 11394 12964 11406
rect 12908 11342 12910 11394
rect 12962 11342 12964 11394
rect 12572 11284 12628 11294
rect 11676 11172 11732 11182
rect 11676 11078 11732 11116
rect 12460 11172 12516 11182
rect 12460 11078 12516 11116
rect 11564 10892 11732 10948
rect 11564 10500 11620 10510
rect 11564 9826 11620 10444
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11564 8036 11620 9774
rect 11676 9266 11732 10892
rect 11900 10500 11956 10510
rect 11900 10406 11956 10444
rect 11676 9214 11678 9266
rect 11730 9214 11732 9266
rect 11676 9202 11732 9214
rect 12124 9828 12180 9838
rect 12124 9714 12180 9772
rect 12124 9662 12126 9714
rect 12178 9662 12180 9714
rect 11564 6802 11620 7980
rect 11564 6750 11566 6802
rect 11618 6750 11620 6802
rect 11564 6738 11620 6750
rect 12012 7588 12068 7598
rect 12012 6580 12068 7532
rect 12124 6692 12180 9662
rect 12236 9156 12292 9166
rect 12236 9062 12292 9100
rect 12572 9044 12628 11228
rect 12796 9940 12852 9950
rect 12684 9716 12740 9726
rect 12684 9622 12740 9660
rect 12796 9714 12852 9884
rect 12796 9662 12798 9714
rect 12850 9662 12852 9714
rect 12796 9380 12852 9662
rect 12796 9314 12852 9324
rect 12684 9044 12740 9054
rect 12572 9042 12740 9044
rect 12572 8990 12686 9042
rect 12738 8990 12740 9042
rect 12572 8988 12740 8990
rect 12684 8372 12740 8988
rect 12908 8596 12964 11342
rect 13020 9604 13076 9614
rect 13020 9510 13076 9548
rect 12908 8530 12964 8540
rect 12796 8372 12852 8382
rect 12684 8370 12852 8372
rect 12684 8318 12798 8370
rect 12850 8318 12852 8370
rect 12684 8316 12852 8318
rect 12796 8306 12852 8316
rect 13132 8260 13188 22092
rect 13692 22148 13748 22158
rect 13692 22146 13860 22148
rect 13692 22094 13694 22146
rect 13746 22094 13860 22146
rect 13692 22092 13860 22094
rect 13692 22082 13748 22092
rect 13244 21474 13300 21486
rect 13244 21422 13246 21474
rect 13298 21422 13300 21474
rect 13244 18564 13300 21422
rect 13692 21474 13748 21486
rect 13692 21422 13694 21474
rect 13746 21422 13748 21474
rect 13580 20580 13636 20590
rect 13692 20580 13748 21422
rect 13804 21026 13860 22092
rect 14028 21810 14084 22204
rect 14700 23042 14756 23054
rect 14700 22990 14702 23042
rect 14754 22990 14756 23042
rect 14140 22148 14196 22158
rect 14140 21924 14196 22092
rect 14140 21858 14196 21868
rect 14028 21758 14030 21810
rect 14082 21758 14084 21810
rect 14028 21746 14084 21758
rect 14700 21588 14756 22990
rect 15148 23042 15204 23054
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 15148 22260 15204 22990
rect 15148 22194 15204 22204
rect 15484 23042 15540 23054
rect 15484 22990 15486 23042
rect 15538 22990 15540 23042
rect 14700 21522 14756 21532
rect 14924 22146 14980 22158
rect 14924 22094 14926 22146
rect 14978 22094 14980 22146
rect 14924 21700 14980 22094
rect 15372 22148 15428 22158
rect 15372 22054 15428 22092
rect 15484 21924 15540 22990
rect 15484 21858 15540 21868
rect 13804 20974 13806 21026
rect 13858 20974 13860 21026
rect 13804 20962 13860 20974
rect 14476 21474 14532 21486
rect 14476 21422 14478 21474
rect 14530 21422 14532 21474
rect 14476 21252 14532 21422
rect 14476 21028 14532 21196
rect 14924 21474 14980 21644
rect 14924 21422 14926 21474
rect 14978 21422 14980 21474
rect 14476 20962 14532 20972
rect 14588 21026 14644 21038
rect 14588 20974 14590 21026
rect 14642 20974 14644 21026
rect 14140 20580 14196 20590
rect 13468 20578 13748 20580
rect 13468 20526 13582 20578
rect 13634 20526 13748 20578
rect 13468 20524 13748 20526
rect 14028 20578 14196 20580
rect 14028 20526 14142 20578
rect 14194 20526 14196 20578
rect 14028 20524 14196 20526
rect 13356 20132 13412 20142
rect 13356 20038 13412 20076
rect 13244 18498 13300 18508
rect 13468 18452 13524 20524
rect 13580 20514 13636 20524
rect 14028 19908 14084 20524
rect 14140 20514 14196 20524
rect 14588 20578 14644 20974
rect 14924 21028 14980 21422
rect 14924 20962 14980 20972
rect 15372 21476 15428 21486
rect 15596 21476 15652 21486
rect 15036 20580 15092 20590
rect 14588 20526 14590 20578
rect 14642 20526 14644 20578
rect 14028 19814 14084 19852
rect 14476 19906 14532 19918
rect 14476 19854 14478 19906
rect 14530 19854 14532 19906
rect 13580 19460 13636 19470
rect 13580 19346 13636 19404
rect 13580 19294 13582 19346
rect 13634 19294 13636 19346
rect 13580 19282 13636 19294
rect 14252 19460 14308 19470
rect 14140 19012 14196 19022
rect 14140 18918 14196 18956
rect 14252 18676 14308 19404
rect 14252 18610 14308 18620
rect 13468 18386 13524 18396
rect 14028 18564 14084 18574
rect 13580 18340 13636 18350
rect 13580 18338 13972 18340
rect 13580 18286 13582 18338
rect 13634 18286 13972 18338
rect 13580 18284 13972 18286
rect 13580 18274 13636 18284
rect 13468 18226 13524 18238
rect 13468 18174 13470 18226
rect 13522 18174 13524 18226
rect 13356 17780 13412 17790
rect 13356 15540 13412 17724
rect 13468 15988 13524 18174
rect 13804 17444 13860 17454
rect 13804 17350 13860 17388
rect 13580 17108 13636 17146
rect 13580 17042 13636 17052
rect 13804 16994 13860 17006
rect 13804 16942 13806 16994
rect 13858 16942 13860 16994
rect 13692 16884 13748 16894
rect 13692 16770 13748 16828
rect 13692 16718 13694 16770
rect 13746 16718 13748 16770
rect 13692 16706 13748 16718
rect 13804 16324 13860 16942
rect 13804 16258 13860 16268
rect 13916 16210 13972 18284
rect 14028 17554 14084 18508
rect 14140 18338 14196 18350
rect 14140 18286 14142 18338
rect 14194 18286 14196 18338
rect 14140 17780 14196 18286
rect 14140 17714 14196 17724
rect 14252 18226 14308 18238
rect 14252 18174 14254 18226
rect 14306 18174 14308 18226
rect 14028 17502 14030 17554
rect 14082 17502 14084 17554
rect 14028 17220 14084 17502
rect 14140 17554 14196 17566
rect 14140 17502 14142 17554
rect 14194 17502 14196 17554
rect 14140 17332 14196 17502
rect 14140 17266 14196 17276
rect 14028 17154 14084 17164
rect 14252 17108 14308 18174
rect 14476 17668 14532 19854
rect 14588 19012 14644 20526
rect 14924 20578 15092 20580
rect 14924 20526 15038 20578
rect 15090 20526 15092 20578
rect 14924 20524 15092 20526
rect 14924 19236 14980 20524
rect 15036 20514 15092 20524
rect 15036 20132 15092 20142
rect 15036 20038 15092 20076
rect 14924 19180 15092 19236
rect 14588 18946 14644 18956
rect 14700 19012 14756 19022
rect 14924 19012 14980 19022
rect 14700 19010 14868 19012
rect 14700 18958 14702 19010
rect 14754 18958 14868 19010
rect 14700 18956 14868 18958
rect 14700 18946 14756 18956
rect 14700 18564 14756 18574
rect 14588 18452 14644 18462
rect 14588 18226 14644 18396
rect 14700 18450 14756 18508
rect 14700 18398 14702 18450
rect 14754 18398 14756 18450
rect 14700 18386 14756 18398
rect 14812 18340 14868 18956
rect 14812 18274 14868 18284
rect 14588 18174 14590 18226
rect 14642 18174 14644 18226
rect 14588 17668 14644 18174
rect 14700 17668 14756 17678
rect 14588 17666 14756 17668
rect 14588 17614 14702 17666
rect 14754 17614 14756 17666
rect 14588 17612 14756 17614
rect 14476 17444 14532 17612
rect 14700 17602 14756 17612
rect 14476 17378 14532 17388
rect 14812 17444 14868 17454
rect 14924 17444 14980 18956
rect 15036 18564 15092 19180
rect 15148 19012 15204 19022
rect 15148 19010 15316 19012
rect 15148 18958 15150 19010
rect 15202 18958 15316 19010
rect 15148 18956 15316 18958
rect 15148 18946 15204 18956
rect 15036 18498 15092 18508
rect 15148 18340 15204 18350
rect 15036 18338 15204 18340
rect 15036 18286 15150 18338
rect 15202 18286 15204 18338
rect 15036 18284 15204 18286
rect 15036 18226 15092 18284
rect 15148 18274 15204 18284
rect 15036 18174 15038 18226
rect 15090 18174 15092 18226
rect 15036 18162 15092 18174
rect 15148 18004 15204 18014
rect 14812 17442 14980 17444
rect 14812 17390 14814 17442
rect 14866 17390 14980 17442
rect 14812 17388 14980 17390
rect 14812 17378 14868 17388
rect 14252 17042 14308 17052
rect 14476 17220 14532 17230
rect 14924 17220 14980 17388
rect 15036 17444 15092 17454
rect 15148 17444 15204 17948
rect 15036 17442 15204 17444
rect 15036 17390 15038 17442
rect 15090 17390 15204 17442
rect 15036 17388 15204 17390
rect 15036 17378 15092 17388
rect 14924 17164 15092 17220
rect 13916 16158 13918 16210
rect 13970 16158 13972 16210
rect 13916 16146 13972 16158
rect 14028 16996 14084 17006
rect 13468 15922 13524 15932
rect 13692 16100 13748 16110
rect 13356 15426 13412 15484
rect 13580 15540 13636 15550
rect 13692 15540 13748 16044
rect 13580 15538 13748 15540
rect 13580 15486 13582 15538
rect 13634 15486 13748 15538
rect 13580 15484 13748 15486
rect 13804 15988 13860 15998
rect 13580 15474 13636 15484
rect 13356 15374 13358 15426
rect 13410 15374 13412 15426
rect 13356 15362 13412 15374
rect 13692 15316 13748 15326
rect 13692 15202 13748 15260
rect 13692 15150 13694 15202
rect 13746 15150 13748 15202
rect 13692 15138 13748 15150
rect 13468 15092 13524 15102
rect 13468 14644 13524 15036
rect 13468 14578 13524 14588
rect 13244 14196 13300 14206
rect 13804 14196 13860 15932
rect 13916 15876 13972 15886
rect 13916 15782 13972 15820
rect 14028 15148 14084 16940
rect 14252 16882 14308 16894
rect 14252 16830 14254 16882
rect 14306 16830 14308 16882
rect 14252 16660 14308 16830
rect 14252 16594 14308 16604
rect 14140 16548 14196 16558
rect 14140 15538 14196 16492
rect 14476 16548 14532 17164
rect 14588 17108 14644 17118
rect 14588 16882 14644 17052
rect 14588 16830 14590 16882
rect 14642 16830 14644 16882
rect 14588 16818 14644 16830
rect 14700 16884 14756 16894
rect 14476 16482 14532 16492
rect 14700 16212 14756 16828
rect 14812 16882 14868 16894
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16660 14868 16830
rect 14812 16594 14868 16604
rect 14924 16882 14980 16894
rect 14924 16830 14926 16882
rect 14978 16830 14980 16882
rect 14924 16324 14980 16830
rect 14924 16258 14980 16268
rect 14140 15486 14142 15538
rect 14194 15486 14196 15538
rect 14140 15474 14196 15486
rect 14476 16156 14756 16212
rect 14028 15092 14308 15148
rect 14140 14644 14196 14654
rect 14028 14532 14084 14542
rect 13244 13858 13300 14140
rect 13468 14140 13860 14196
rect 13916 14476 14028 14532
rect 13244 13806 13246 13858
rect 13298 13806 13300 13858
rect 13244 13794 13300 13806
rect 13356 13858 13412 13870
rect 13356 13806 13358 13858
rect 13410 13806 13412 13858
rect 13356 13748 13412 13806
rect 13356 13682 13412 13692
rect 13468 11508 13524 14140
rect 13580 13972 13636 13982
rect 13916 13972 13972 14476
rect 14028 14438 14084 14476
rect 14140 14418 14196 14588
rect 14140 14366 14142 14418
rect 14194 14366 14196 14418
rect 14140 14354 14196 14366
rect 13580 13970 13972 13972
rect 13580 13918 13582 13970
rect 13634 13918 13972 13970
rect 13580 13916 13972 13918
rect 13580 13906 13636 13916
rect 14252 13076 14308 15092
rect 14476 14980 14532 16156
rect 14588 15988 14644 15998
rect 14588 15894 14644 15932
rect 14700 15986 14756 16156
rect 14700 15934 14702 15986
rect 14754 15934 14756 15986
rect 14700 15922 14756 15934
rect 14812 16100 14868 16110
rect 14812 15764 14868 16044
rect 14812 15698 14868 15708
rect 14924 15988 14980 15998
rect 14924 15874 14980 15932
rect 14924 15822 14926 15874
rect 14978 15822 14980 15874
rect 14588 15652 14644 15662
rect 14588 15316 14644 15596
rect 14588 15250 14644 15260
rect 14700 15540 14756 15550
rect 14700 15148 14756 15484
rect 14924 15314 14980 15822
rect 14924 15262 14926 15314
rect 14978 15262 14980 15314
rect 14924 15250 14980 15262
rect 14476 14914 14532 14924
rect 14588 15092 14756 15148
rect 14812 15202 14868 15214
rect 14812 15150 14814 15202
rect 14866 15150 14868 15202
rect 14588 14420 14644 15092
rect 14812 14644 14868 15150
rect 15036 14756 15092 17164
rect 15260 17108 15316 18956
rect 15372 17892 15428 21420
rect 15484 21474 15652 21476
rect 15484 21422 15598 21474
rect 15650 21422 15652 21474
rect 15484 21420 15652 21422
rect 15484 19572 15540 21420
rect 15596 21410 15652 21420
rect 15820 20578 15876 20590
rect 15820 20526 15822 20578
rect 15874 20526 15876 20578
rect 15596 19908 15652 19918
rect 15596 19906 15764 19908
rect 15596 19854 15598 19906
rect 15650 19854 15764 19906
rect 15596 19852 15764 19854
rect 15596 19842 15652 19852
rect 15484 19506 15540 19516
rect 15596 19012 15652 19022
rect 15372 17826 15428 17836
rect 15484 19010 15652 19012
rect 15484 18958 15598 19010
rect 15650 18958 15652 19010
rect 15484 18956 15652 18958
rect 15484 18226 15540 18956
rect 15596 18946 15652 18956
rect 15708 18676 15764 19852
rect 15708 18610 15764 18620
rect 15484 18174 15486 18226
rect 15538 18174 15540 18226
rect 15148 17052 15316 17108
rect 15372 17668 15428 17678
rect 15148 15764 15204 17052
rect 15372 16996 15428 17612
rect 15372 16930 15428 16940
rect 15260 16882 15316 16894
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16772 15316 16830
rect 15260 16706 15316 16716
rect 15372 16770 15428 16782
rect 15372 16718 15374 16770
rect 15426 16718 15428 16770
rect 15372 16548 15428 16718
rect 15484 16660 15540 18174
rect 15596 18340 15652 18350
rect 15596 16884 15652 18284
rect 15820 18228 15876 20526
rect 15932 20132 15988 32284
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 20972 25284 21028 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19516 24276 19572 24286
rect 19404 24052 19460 24062
rect 17612 23828 17668 23838
rect 16828 23156 16884 23166
rect 16828 23062 16884 23100
rect 16044 23042 16100 23054
rect 16044 22990 16046 23042
rect 16098 22990 16100 23042
rect 16044 22372 16100 22990
rect 16492 23042 16548 23054
rect 16492 22990 16494 23042
rect 16546 22990 16548 23042
rect 16492 22820 16548 22990
rect 16940 23044 16996 23054
rect 16492 22754 16548 22764
rect 16828 22820 16884 22830
rect 16044 22306 16100 22316
rect 16492 22260 16548 22270
rect 16492 22166 16548 22204
rect 16156 22148 16212 22158
rect 16156 21924 16212 22092
rect 16156 21858 16212 21868
rect 16828 21812 16884 22764
rect 16940 22148 16996 22988
rect 17388 22484 17444 22494
rect 17388 22390 17444 22428
rect 16940 22054 16996 22092
rect 16940 21812 16996 21822
rect 16828 21810 16996 21812
rect 16828 21758 16942 21810
rect 16994 21758 16996 21810
rect 16828 21756 16996 21758
rect 16940 21746 16996 21756
rect 17612 21812 17668 23772
rect 17836 22596 17892 22606
rect 17836 22482 17892 22540
rect 17836 22430 17838 22482
rect 17890 22430 17892 22482
rect 17836 22418 17892 22430
rect 16044 21700 16100 21710
rect 16044 21606 16100 21644
rect 16492 21700 16548 21710
rect 17612 21680 17668 21756
rect 18060 22260 18116 22270
rect 16492 21606 16548 21644
rect 15932 20066 15988 20076
rect 16156 21588 16212 21598
rect 16156 20356 16212 21532
rect 16268 20580 16324 20590
rect 16268 20486 16324 20524
rect 16604 20578 16660 20590
rect 16604 20526 16606 20578
rect 16658 20526 16660 20578
rect 16044 19906 16100 19918
rect 16044 19854 16046 19906
rect 16098 19854 16100 19906
rect 15820 18162 15876 18172
rect 15932 19010 15988 19022
rect 15932 18958 15934 19010
rect 15986 18958 15988 19010
rect 15932 18788 15988 18958
rect 16044 19012 16100 19854
rect 16044 18946 16100 18956
rect 16156 18788 16212 20300
rect 16604 20244 16660 20526
rect 16604 20178 16660 20188
rect 16940 20580 16996 20590
rect 16716 19908 16772 19918
rect 16716 19814 16772 19852
rect 16940 19796 16996 20524
rect 17388 20578 17444 20590
rect 17388 20526 17390 20578
rect 17442 20526 17444 20578
rect 17388 20356 17444 20526
rect 17948 20580 18004 20590
rect 17948 20486 18004 20524
rect 17388 20290 17444 20300
rect 15932 18732 16212 18788
rect 16380 19012 16436 19022
rect 15596 16818 15652 16828
rect 15708 18004 15764 18014
rect 15708 16882 15764 17948
rect 15932 17220 15988 18732
rect 16156 18338 16212 18350
rect 16156 18286 16158 18338
rect 16210 18286 16212 18338
rect 16156 18004 16212 18286
rect 16156 17938 16212 17948
rect 15932 17154 15988 17164
rect 16044 17442 16100 17454
rect 16044 17390 16046 17442
rect 16098 17390 16100 17442
rect 16044 16996 16100 17390
rect 16044 16930 16100 16940
rect 16156 17108 16212 17118
rect 15708 16830 15710 16882
rect 15762 16830 15764 16882
rect 15708 16818 15764 16830
rect 15820 16882 15876 16894
rect 15820 16830 15822 16882
rect 15874 16830 15876 16882
rect 15484 16604 15652 16660
rect 15148 15698 15204 15708
rect 15260 16492 15428 16548
rect 15260 15540 15316 16492
rect 15372 15988 15428 15998
rect 15372 15894 15428 15932
rect 15036 14690 15092 14700
rect 15148 15484 15316 15540
rect 14812 14512 14868 14588
rect 15036 14532 15092 14542
rect 15036 14438 15092 14476
rect 14364 14306 14420 14318
rect 14364 14254 14366 14306
rect 14418 14254 14420 14306
rect 14364 13858 14420 14254
rect 14588 13970 14644 14364
rect 14588 13918 14590 13970
rect 14642 13918 14644 13970
rect 14588 13906 14644 13918
rect 15148 13972 15204 15484
rect 15260 15316 15316 15354
rect 15260 15250 15316 15260
rect 15372 14306 15428 14318
rect 15372 14254 15374 14306
rect 15426 14254 15428 14306
rect 15148 13906 15204 13916
rect 15260 14196 15316 14206
rect 14364 13806 14366 13858
rect 14418 13806 14420 13858
rect 14364 13794 14420 13806
rect 14812 13858 14868 13870
rect 14812 13806 14814 13858
rect 14866 13806 14868 13858
rect 14476 13524 14532 13534
rect 14476 13430 14532 13468
rect 14812 13524 14868 13806
rect 14812 13458 14868 13468
rect 14924 13636 14980 13646
rect 14364 13188 14420 13198
rect 14364 13094 14420 13132
rect 14924 13186 14980 13580
rect 14924 13134 14926 13186
rect 14978 13134 14980 13186
rect 14924 13122 14980 13134
rect 15036 13300 15092 13310
rect 14028 13020 14308 13076
rect 14588 13076 14644 13086
rect 13692 12852 13748 12862
rect 13692 12758 13748 12796
rect 13468 11452 13860 11508
rect 13692 11282 13748 11294
rect 13692 11230 13694 11282
rect 13746 11230 13748 11282
rect 13356 10052 13412 10062
rect 13692 10052 13748 11230
rect 13412 9996 13748 10052
rect 13356 9154 13412 9996
rect 13692 9828 13748 9838
rect 13804 9828 13860 11452
rect 14028 11506 14084 13020
rect 14588 12962 14644 13020
rect 14588 12910 14590 12962
rect 14642 12910 14644 12962
rect 14028 11454 14030 11506
rect 14082 11454 14084 11506
rect 14028 11172 14084 11454
rect 14028 11106 14084 11116
rect 14252 12850 14308 12862
rect 14252 12798 14254 12850
rect 14306 12798 14308 12850
rect 14028 10498 14084 10510
rect 14028 10446 14030 10498
rect 14082 10446 14084 10498
rect 14028 9938 14084 10446
rect 14252 10164 14308 12798
rect 14588 12404 14644 12910
rect 14812 12964 14868 12974
rect 14812 12870 14868 12908
rect 14588 12338 14644 12348
rect 14588 12068 14644 12078
rect 14588 10612 14644 12012
rect 14924 11620 14980 11630
rect 14700 11284 14756 11294
rect 14700 11190 14756 11228
rect 14812 11170 14868 11182
rect 14812 11118 14814 11170
rect 14866 11118 14868 11170
rect 14812 10836 14868 11118
rect 14700 10612 14756 10622
rect 14588 10610 14756 10612
rect 14588 10558 14702 10610
rect 14754 10558 14756 10610
rect 14588 10556 14756 10558
rect 14700 10546 14756 10556
rect 14812 10276 14868 10780
rect 14252 10098 14308 10108
rect 14588 10220 14868 10276
rect 14924 10500 14980 11564
rect 14028 9886 14030 9938
rect 14082 9886 14084 9938
rect 14028 9874 14084 9886
rect 14140 10052 14196 10062
rect 13916 9828 13972 9838
rect 13804 9772 13916 9828
rect 13468 9268 13524 9278
rect 13468 9174 13524 9212
rect 13356 9102 13358 9154
rect 13410 9102 13412 9154
rect 13356 9090 13412 9102
rect 12684 7700 12740 7710
rect 12348 6804 12404 6814
rect 12236 6692 12292 6702
rect 12124 6690 12292 6692
rect 12124 6638 12238 6690
rect 12290 6638 12292 6690
rect 12124 6636 12292 6638
rect 12236 6626 12292 6636
rect 12012 6524 12180 6580
rect 11564 6020 11620 6030
rect 11564 5926 11620 5964
rect 10556 4286 10558 4338
rect 10610 4286 10612 4338
rect 10556 4274 10612 4286
rect 10108 3726 10110 3778
rect 10162 3726 10164 3778
rect 10108 3714 10164 3726
rect 10332 4228 10388 4238
rect 10332 3778 10388 4172
rect 11228 4226 11284 4238
rect 11228 4174 11230 4226
rect 11282 4174 11284 4226
rect 11228 4116 11284 4174
rect 11228 4050 11284 4060
rect 10668 3892 10724 3902
rect 10332 3726 10334 3778
rect 10386 3726 10388 3778
rect 10332 3714 10388 3726
rect 10556 3780 10612 3790
rect 10556 3686 10612 3724
rect 10668 3778 10724 3836
rect 11452 3892 11508 5740
rect 11900 5460 11956 5470
rect 11900 5010 11956 5404
rect 11900 4958 11902 5010
rect 11954 4958 11956 5010
rect 11900 4946 11956 4958
rect 12012 5346 12068 5358
rect 12012 5294 12014 5346
rect 12066 5294 12068 5346
rect 12012 4564 12068 5294
rect 12124 5010 12180 6524
rect 12348 6020 12404 6748
rect 12684 6690 12740 7644
rect 13132 7586 13188 8204
rect 13580 8932 13636 8942
rect 13580 7924 13636 8876
rect 13692 8372 13748 9772
rect 13916 9696 13972 9772
rect 14140 9826 14196 9996
rect 14140 9774 14142 9826
rect 14194 9774 14196 9826
rect 14140 9762 14196 9774
rect 14252 9940 14308 9950
rect 14252 9268 14308 9884
rect 14364 9828 14420 9838
rect 14364 9826 14532 9828
rect 14364 9774 14366 9826
rect 14418 9774 14532 9826
rect 14364 9772 14532 9774
rect 14364 9762 14420 9772
rect 14028 9212 14420 9268
rect 14028 9154 14084 9212
rect 14028 9102 14030 9154
rect 14082 9102 14084 9154
rect 14028 9090 14084 9102
rect 14252 9042 14308 9054
rect 14252 8990 14254 9042
rect 14306 8990 14308 9042
rect 13804 8820 13860 8830
rect 13804 8818 13972 8820
rect 13804 8766 13806 8818
rect 13858 8766 13972 8818
rect 13804 8764 13972 8766
rect 13804 8754 13860 8764
rect 13692 8306 13748 8316
rect 13804 8596 13860 8606
rect 13804 8370 13860 8540
rect 13916 8484 13972 8764
rect 14140 8484 14196 8494
rect 13916 8482 14196 8484
rect 13916 8430 14142 8482
rect 14194 8430 14196 8482
rect 13916 8428 14196 8430
rect 13804 8318 13806 8370
rect 13858 8318 13860 8370
rect 13804 8306 13860 8318
rect 13916 8258 13972 8270
rect 13916 8206 13918 8258
rect 13970 8206 13972 8258
rect 13692 8148 13748 8158
rect 13692 8054 13748 8092
rect 13916 7924 13972 8206
rect 14140 8260 14196 8428
rect 14140 8036 14196 8204
rect 14140 7970 14196 7980
rect 13580 7868 13972 7924
rect 13132 7534 13134 7586
rect 13186 7534 13188 7586
rect 13132 7522 13188 7534
rect 12684 6638 12686 6690
rect 12738 6638 12740 6690
rect 12684 6626 12740 6638
rect 13804 6692 13860 6702
rect 12460 6580 12516 6590
rect 12460 6486 12516 6524
rect 13804 6578 13860 6636
rect 13804 6526 13806 6578
rect 13858 6526 13860 6578
rect 13804 6514 13860 6526
rect 12572 6468 12628 6478
rect 12796 6468 12852 6478
rect 12572 6466 12740 6468
rect 12572 6414 12574 6466
rect 12626 6414 12740 6466
rect 12572 6412 12740 6414
rect 12572 6402 12628 6412
rect 12124 4958 12126 5010
rect 12178 4958 12180 5010
rect 12124 4946 12180 4958
rect 12236 6018 12404 6020
rect 12236 5966 12350 6018
rect 12402 5966 12404 6018
rect 12236 5964 12404 5966
rect 12012 4498 12068 4508
rect 11452 3826 11508 3836
rect 10668 3726 10670 3778
rect 10722 3726 10724 3778
rect 10668 3714 10724 3726
rect 11676 3556 11732 3566
rect 11676 3442 11732 3500
rect 11676 3390 11678 3442
rect 11730 3390 11732 3442
rect 11676 3378 11732 3390
rect 12236 3388 12292 5964
rect 12348 5954 12404 5964
rect 12572 5124 12628 5134
rect 12572 5030 12628 5068
rect 12348 5012 12404 5022
rect 12348 4918 12404 4956
rect 12684 4340 12740 6412
rect 12796 6374 12852 6412
rect 13916 6356 13972 7868
rect 14140 6580 14196 6590
rect 14140 6486 14196 6524
rect 13916 6290 13972 6300
rect 14252 6020 14308 8990
rect 14364 8258 14420 9212
rect 14364 8206 14366 8258
rect 14418 8206 14420 8258
rect 14364 6690 14420 8206
rect 14476 7812 14532 9772
rect 14476 7746 14532 7756
rect 14588 9492 14644 10220
rect 14924 10164 14980 10444
rect 14364 6638 14366 6690
rect 14418 6638 14420 6690
rect 14364 6244 14420 6638
rect 14588 6580 14644 9436
rect 14812 10108 14980 10164
rect 14812 9716 14868 10108
rect 15036 10052 15092 13244
rect 14924 9996 15092 10052
rect 14924 9940 14980 9996
rect 14924 9874 14980 9884
rect 15036 9828 15092 9838
rect 14924 9716 14980 9726
rect 14812 9714 14980 9716
rect 14812 9662 14926 9714
rect 14978 9662 14980 9714
rect 14812 9660 14980 9662
rect 14700 9380 14756 9390
rect 14700 9266 14756 9324
rect 14700 9214 14702 9266
rect 14754 9214 14756 9266
rect 14700 9202 14756 9214
rect 14588 6514 14644 6524
rect 14700 8258 14756 8270
rect 14700 8206 14702 8258
rect 14754 8206 14756 8258
rect 14364 6178 14420 6188
rect 14028 5964 14308 6020
rect 13468 5796 13524 5806
rect 13468 5702 13524 5740
rect 13692 4900 13748 4910
rect 12684 4274 12740 4284
rect 13356 4898 13748 4900
rect 13356 4846 13694 4898
rect 13746 4846 13748 4898
rect 13356 4844 13748 4846
rect 13356 4226 13412 4844
rect 13692 4834 13748 4844
rect 13916 4452 13972 4462
rect 13916 4338 13972 4396
rect 13916 4286 13918 4338
rect 13970 4286 13972 4338
rect 13916 4274 13972 4286
rect 13356 4174 13358 4226
rect 13410 4174 13412 4226
rect 13356 4162 13412 4174
rect 14028 3778 14084 5964
rect 14140 5794 14196 5806
rect 14700 5796 14756 8206
rect 14812 8148 14868 9660
rect 14924 9650 14980 9660
rect 15036 9602 15092 9772
rect 15260 9828 15316 14140
rect 15372 13858 15428 14254
rect 15372 13806 15374 13858
rect 15426 13806 15428 13858
rect 15372 13524 15428 13806
rect 15596 13748 15652 16604
rect 15820 16100 15876 16830
rect 16156 16212 16212 17052
rect 16268 16884 16324 16894
rect 16268 16790 16324 16828
rect 16380 16324 16436 18956
rect 16604 19012 16660 19022
rect 16604 19010 16772 19012
rect 16604 18958 16606 19010
rect 16658 18958 16772 19010
rect 16604 18956 16772 18958
rect 16604 18946 16660 18956
rect 16604 18338 16660 18350
rect 16604 18286 16606 18338
rect 16658 18286 16660 18338
rect 16604 18226 16660 18286
rect 16604 18174 16606 18226
rect 16658 18174 16660 18226
rect 16604 18162 16660 18174
rect 16492 17892 16548 17902
rect 16492 17108 16548 17836
rect 16492 16976 16548 17052
rect 16604 16884 16660 16894
rect 16716 16884 16772 18956
rect 16940 19010 16996 19740
rect 17612 19908 17668 19918
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 16940 18900 16996 18958
rect 17388 19012 17444 19022
rect 17388 18918 17444 18956
rect 16940 18834 16996 18844
rect 17052 18564 17108 18574
rect 16828 17892 16884 17902
rect 16828 17778 16884 17836
rect 16828 17726 16830 17778
rect 16882 17726 16884 17778
rect 16828 17714 16884 17726
rect 16660 16828 16772 16884
rect 16940 16996 16996 17006
rect 16604 16790 16660 16828
rect 16380 16268 16772 16324
rect 16156 16156 16660 16212
rect 15708 15988 15764 15998
rect 15708 15894 15764 15932
rect 15708 15764 15764 15774
rect 15708 15314 15764 15708
rect 15708 15262 15710 15314
rect 15762 15262 15764 15314
rect 15708 15250 15764 15262
rect 15820 15204 15876 16044
rect 16492 15986 16548 15998
rect 16492 15934 16494 15986
rect 16546 15934 16548 15986
rect 16156 15876 16212 15886
rect 16156 15874 16324 15876
rect 16156 15822 16158 15874
rect 16210 15822 16324 15874
rect 16156 15820 16324 15822
rect 16156 15810 16212 15820
rect 16156 15314 16212 15326
rect 16156 15262 16158 15314
rect 16210 15262 16212 15314
rect 15820 15138 15876 15148
rect 15932 15202 15988 15214
rect 15932 15150 15934 15202
rect 15986 15150 15988 15202
rect 15932 14644 15988 15150
rect 16156 15204 16212 15262
rect 16268 15314 16324 15820
rect 16380 15874 16436 15886
rect 16380 15822 16382 15874
rect 16434 15822 16436 15874
rect 16380 15764 16436 15822
rect 16380 15698 16436 15708
rect 16492 15540 16548 15934
rect 16268 15262 16270 15314
rect 16322 15262 16324 15314
rect 16268 15250 16324 15262
rect 16380 15484 16492 15540
rect 16156 15138 16212 15148
rect 16268 14756 16324 14766
rect 16380 14756 16436 15484
rect 16492 15474 16548 15484
rect 16268 14754 16436 14756
rect 16268 14702 16270 14754
rect 16322 14702 16436 14754
rect 16268 14700 16436 14702
rect 16268 14690 16324 14700
rect 15932 14578 15988 14588
rect 16268 14532 16324 14542
rect 16268 14438 16324 14476
rect 15932 14420 15988 14430
rect 16604 14420 16660 16156
rect 15372 13458 15428 13468
rect 15484 13634 15540 13646
rect 15484 13582 15486 13634
rect 15538 13582 15540 13634
rect 15372 11620 15428 11630
rect 15372 10836 15428 11564
rect 15372 10722 15428 10780
rect 15484 10834 15540 13582
rect 15596 12628 15652 13692
rect 15708 14418 15988 14420
rect 15708 14366 15934 14418
rect 15986 14366 15988 14418
rect 15708 14364 15988 14366
rect 15708 13860 15764 14364
rect 15932 14354 15988 14364
rect 16380 14364 16660 14420
rect 16380 14308 16436 14364
rect 16268 14252 16436 14308
rect 15820 13860 15876 13870
rect 15708 13804 15820 13860
rect 15708 12962 15764 13804
rect 15820 13766 15876 13804
rect 15708 12910 15710 12962
rect 15762 12910 15764 12962
rect 15708 12898 15764 12910
rect 15820 13524 15876 13534
rect 15820 12962 15876 13468
rect 16268 13188 16324 14252
rect 16716 14196 16772 16268
rect 16828 15540 16884 15550
rect 16828 14530 16884 15484
rect 16940 15538 16996 16940
rect 16940 15486 16942 15538
rect 16994 15486 16996 15538
rect 16940 15474 16996 15486
rect 17052 15148 17108 18508
rect 17612 18564 17668 19852
rect 17948 19906 18004 19918
rect 17948 19854 17950 19906
rect 18002 19854 18004 19906
rect 17836 19348 17892 19358
rect 17948 19348 18004 19854
rect 17892 19292 18004 19348
rect 17836 19282 17892 19292
rect 17612 18450 17668 18508
rect 17612 18398 17614 18450
rect 17666 18398 17668 18450
rect 17612 18386 17668 18398
rect 17388 18228 17444 18238
rect 17388 17778 17444 18172
rect 17948 18116 18004 19292
rect 18060 19348 18116 22204
rect 18284 22148 18340 22158
rect 18284 22054 18340 22092
rect 18284 21924 18340 21934
rect 18172 21476 18228 21486
rect 18172 21382 18228 21420
rect 18284 20578 18340 21868
rect 19404 21810 19460 23996
rect 19404 21758 19406 21810
rect 19458 21758 19460 21810
rect 19404 21746 19460 21758
rect 18508 21476 18564 21486
rect 18508 21382 18564 21420
rect 18956 21474 19012 21486
rect 18956 21422 18958 21474
rect 19010 21422 19012 21474
rect 18284 20526 18286 20578
rect 18338 20526 18340 20578
rect 18284 20242 18340 20526
rect 18732 20580 18788 20590
rect 18732 20486 18788 20524
rect 18284 20190 18286 20242
rect 18338 20190 18340 20242
rect 18284 20178 18340 20190
rect 18956 20188 19012 21422
rect 19180 20578 19236 20590
rect 19180 20526 19182 20578
rect 19234 20526 19236 20578
rect 18060 19216 18116 19292
rect 18172 20132 18228 20142
rect 18956 20132 19124 20188
rect 17388 17726 17390 17778
rect 17442 17726 17444 17778
rect 17388 16996 17444 17726
rect 17388 16930 17444 16940
rect 17612 18060 18004 18116
rect 18060 18676 18116 18686
rect 17612 16212 17668 18060
rect 18060 17780 18116 18620
rect 18172 18452 18228 20076
rect 18732 19908 18788 19918
rect 18508 19906 18788 19908
rect 18508 19854 18734 19906
rect 18786 19854 18788 19906
rect 18508 19852 18788 19854
rect 18508 19124 18564 19852
rect 18732 19842 18788 19852
rect 18508 19030 18564 19068
rect 18620 19572 18676 19582
rect 18172 18320 18228 18396
rect 18620 18338 18676 19516
rect 18956 19124 19012 19134
rect 18956 19030 19012 19068
rect 18620 18286 18622 18338
rect 18674 18286 18676 18338
rect 18060 17778 18228 17780
rect 18060 17726 18062 17778
rect 18114 17726 18228 17778
rect 18060 17724 18228 17726
rect 18060 17714 18116 17724
rect 18172 17444 18228 17724
rect 18172 17388 18452 17444
rect 17724 16996 17780 17006
rect 17724 16436 17780 16940
rect 18396 16994 18452 17388
rect 18508 17442 18564 17454
rect 18508 17390 18510 17442
rect 18562 17390 18564 17442
rect 18508 17220 18564 17390
rect 18508 17154 18564 17164
rect 18396 16942 18398 16994
rect 18450 16942 18452 16994
rect 18396 16930 18452 16942
rect 18508 16996 18564 17006
rect 18508 16902 18564 16940
rect 17836 16660 17892 16670
rect 17836 16658 18228 16660
rect 17836 16606 17838 16658
rect 17890 16606 18228 16658
rect 17836 16604 18228 16606
rect 17836 16594 17892 16604
rect 17724 16380 18116 16436
rect 17612 16156 17780 16212
rect 17164 15988 17220 15998
rect 17164 15894 17220 15932
rect 17388 15986 17444 15998
rect 17388 15934 17390 15986
rect 17442 15934 17444 15986
rect 17276 15874 17332 15886
rect 17276 15822 17278 15874
rect 17330 15822 17332 15874
rect 16828 14478 16830 14530
rect 16882 14478 16884 14530
rect 16828 14466 16884 14478
rect 16940 15092 17108 15148
rect 17164 15652 17220 15662
rect 16716 14130 16772 14140
rect 16604 13972 16660 13982
rect 16268 13132 16436 13188
rect 15820 12910 15822 12962
rect 15874 12910 15876 12962
rect 15820 12898 15876 12910
rect 16268 12962 16324 12974
rect 16268 12910 16270 12962
rect 16322 12910 16324 12962
rect 15596 12562 15652 12572
rect 15932 12738 15988 12750
rect 15932 12686 15934 12738
rect 15986 12686 15988 12738
rect 15820 12516 15876 12526
rect 15708 11284 15764 11294
rect 15484 10782 15486 10834
rect 15538 10782 15540 10834
rect 15484 10770 15540 10782
rect 15596 11170 15652 11182
rect 15596 11118 15598 11170
rect 15650 11118 15652 11170
rect 15372 10670 15374 10722
rect 15426 10670 15428 10722
rect 15372 10658 15428 10670
rect 15596 10052 15652 11118
rect 15708 10834 15764 11228
rect 15820 10948 15876 12460
rect 15932 11618 15988 12686
rect 16268 12628 16324 12910
rect 16268 12562 16324 12572
rect 15932 11566 15934 11618
rect 15986 11566 15988 11618
rect 15932 11554 15988 11566
rect 16268 12292 16324 12302
rect 16268 11396 16324 12236
rect 16156 11284 16212 11294
rect 16156 11190 16212 11228
rect 15820 10882 15876 10892
rect 15708 10782 15710 10834
rect 15762 10782 15764 10834
rect 15708 10770 15764 10782
rect 16156 10836 16212 10846
rect 15596 9986 15652 9996
rect 16044 9940 16100 9950
rect 16044 9846 16100 9884
rect 15260 9762 15316 9772
rect 16156 9826 16212 10780
rect 16268 10834 16324 11340
rect 16268 10782 16270 10834
rect 16322 10782 16324 10834
rect 16268 10770 16324 10782
rect 16380 10834 16436 13132
rect 16604 12962 16660 13916
rect 16828 13858 16884 13870
rect 16828 13806 16830 13858
rect 16882 13806 16884 13858
rect 16716 13748 16772 13758
rect 16716 13654 16772 13692
rect 16828 13188 16884 13806
rect 16828 13122 16884 13132
rect 16940 12964 16996 15092
rect 17052 14532 17108 14542
rect 17164 14532 17220 15596
rect 17276 15428 17332 15822
rect 17276 15362 17332 15372
rect 17388 14754 17444 15934
rect 17612 15314 17668 15326
rect 17612 15262 17614 15314
rect 17666 15262 17668 15314
rect 17612 15148 17668 15262
rect 17388 14702 17390 14754
rect 17442 14702 17444 14754
rect 17388 14690 17444 14702
rect 17500 15092 17668 15148
rect 17052 14530 17220 14532
rect 17052 14478 17054 14530
rect 17106 14478 17220 14530
rect 17052 14476 17220 14478
rect 17052 14466 17108 14476
rect 17276 14308 17332 14318
rect 17276 14214 17332 14252
rect 17052 14196 17108 14206
rect 17052 13970 17108 14140
rect 17500 13972 17556 15092
rect 17052 13918 17054 13970
rect 17106 13918 17108 13970
rect 17052 13906 17108 13918
rect 17164 13916 17556 13972
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 12898 16660 12910
rect 16716 12908 16996 12964
rect 16716 12180 16772 12908
rect 17164 12850 17220 13916
rect 17164 12798 17166 12850
rect 17218 12798 17220 12850
rect 17164 12786 17220 12798
rect 17388 13188 17444 13198
rect 17388 12850 17444 13132
rect 17724 13076 17780 16156
rect 17948 16100 18004 16110
rect 17948 16006 18004 16044
rect 18060 15986 18116 16380
rect 18060 15934 18062 15986
rect 18114 15934 18116 15986
rect 18060 15922 18116 15934
rect 17836 15540 17892 15550
rect 17836 15446 17892 15484
rect 17948 15316 18004 15326
rect 17948 15222 18004 15260
rect 18172 14532 18228 16604
rect 18284 15876 18340 15886
rect 18620 15876 18676 18286
rect 19068 18452 19124 20132
rect 19180 18564 19236 20526
rect 19516 20132 19572 24220
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21812 20356 21822
rect 19628 20692 19684 20702
rect 19628 20598 19684 20636
rect 20076 20580 20132 20590
rect 20076 20578 20244 20580
rect 20076 20526 20078 20578
rect 20130 20526 20244 20578
rect 20076 20524 20244 20526
rect 20076 20514 20132 20524
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19852 20244 19908 20254
rect 19516 20076 19796 20132
rect 19292 19908 19348 19918
rect 19628 19908 19684 19918
rect 19292 19814 19348 19852
rect 19404 19906 19684 19908
rect 19404 19854 19630 19906
rect 19682 19854 19684 19906
rect 19404 19852 19684 19854
rect 19404 19348 19460 19852
rect 19628 19842 19684 19852
rect 19404 19254 19460 19292
rect 19740 19012 19796 20076
rect 19180 18498 19236 18508
rect 19628 18956 19796 19012
rect 19852 19012 19908 20188
rect 20076 19908 20132 19918
rect 20076 19814 20132 19852
rect 18956 17890 19012 17902
rect 18956 17838 18958 17890
rect 19010 17838 19012 17890
rect 18956 17778 19012 17838
rect 18956 17726 18958 17778
rect 19010 17726 19012 17778
rect 18732 17108 18788 17118
rect 18732 17014 18788 17052
rect 18844 16324 18900 16334
rect 18844 16230 18900 16268
rect 18732 15988 18788 16026
rect 18732 15922 18788 15932
rect 18340 15820 18676 15876
rect 18844 15876 18900 15886
rect 18284 15782 18340 15820
rect 18844 15764 18900 15820
rect 18732 15708 18900 15764
rect 18732 15540 18788 15708
rect 18956 15652 19012 17726
rect 19068 17556 19124 18396
rect 19628 18450 19684 18956
rect 19852 18946 19908 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18676 20244 20524
rect 20300 19348 20356 21756
rect 20524 20916 20580 20926
rect 20524 20242 20580 20860
rect 20524 20190 20526 20242
rect 20578 20190 20580 20242
rect 20524 20178 20580 20190
rect 20972 20130 21028 25228
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 42700 23940 42756 23950
rect 20972 20078 20974 20130
rect 21026 20078 21028 20130
rect 20972 20066 21028 20078
rect 21308 23156 21364 23166
rect 20300 19216 20356 19292
rect 20748 19012 20804 19022
rect 20748 19010 21028 19012
rect 20748 18958 20750 19010
rect 20802 18958 21028 19010
rect 20748 18956 21028 18958
rect 20748 18946 20804 18956
rect 20188 18620 20356 18676
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 19068 17490 19124 17500
rect 19180 18340 19236 18350
rect 19068 16996 19124 17006
rect 19068 16902 19124 16940
rect 18620 15484 18788 15540
rect 18844 15596 19012 15652
rect 19068 15988 19124 15998
rect 18396 15428 18452 15438
rect 18172 14476 18340 14532
rect 18060 14418 18116 14430
rect 18060 14366 18062 14418
rect 18114 14366 18116 14418
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 17388 12786 17444 12798
rect 17500 13020 17780 13076
rect 17836 14308 17892 14318
rect 16940 12738 16996 12750
rect 16940 12686 16942 12738
rect 16994 12686 16996 12738
rect 16940 12628 16996 12686
rect 16940 12562 16996 12572
rect 17276 12738 17332 12750
rect 17276 12686 17278 12738
rect 17330 12686 17332 12738
rect 16604 12178 16772 12180
rect 16604 12126 16718 12178
rect 16770 12126 16772 12178
rect 16604 12124 16772 12126
rect 16380 10782 16382 10834
rect 16434 10782 16436 10834
rect 16380 10612 16436 10782
rect 16492 11172 16548 11182
rect 16492 10722 16548 11116
rect 16492 10670 16494 10722
rect 16546 10670 16548 10722
rect 16492 10658 16548 10670
rect 16380 10546 16436 10556
rect 16604 10500 16660 12124
rect 16716 12114 16772 12124
rect 16940 12404 16996 12414
rect 16156 9774 16158 9826
rect 16210 9774 16212 9826
rect 16156 9762 16212 9774
rect 16268 10388 16324 10398
rect 15036 9550 15038 9602
rect 15090 9550 15092 9602
rect 15036 9538 15092 9550
rect 15148 9492 15204 9502
rect 15148 9044 15204 9436
rect 15260 9268 15316 9278
rect 16156 9268 16212 9278
rect 15260 9266 16212 9268
rect 15260 9214 15262 9266
rect 15314 9214 16158 9266
rect 16210 9214 16212 9266
rect 15260 9212 16212 9214
rect 15260 9202 15316 9212
rect 16156 9202 16212 9212
rect 16268 9266 16324 10332
rect 16268 9214 16270 9266
rect 16322 9214 16324 9266
rect 16268 9202 16324 9214
rect 16492 9828 16548 9838
rect 15484 9044 15540 9054
rect 15148 8988 15316 9044
rect 15148 8820 15204 8830
rect 15148 8370 15204 8764
rect 15260 8482 15316 8988
rect 15260 8430 15262 8482
rect 15314 8430 15316 8482
rect 15260 8418 15316 8430
rect 15372 8930 15428 8942
rect 15372 8878 15374 8930
rect 15426 8878 15428 8930
rect 15148 8318 15150 8370
rect 15202 8318 15204 8370
rect 15148 8306 15204 8318
rect 14812 8082 14868 8092
rect 15260 7812 15316 7822
rect 15260 6802 15316 7756
rect 15372 7700 15428 8878
rect 15484 8596 15540 8988
rect 15820 9044 15876 9054
rect 15820 8950 15876 8988
rect 16492 9044 16548 9772
rect 16492 8950 16548 8988
rect 15484 8530 15540 8540
rect 15820 8484 15876 8494
rect 15820 8370 15876 8428
rect 15820 8318 15822 8370
rect 15874 8318 15876 8370
rect 15820 8306 15876 8318
rect 15372 7634 15428 7644
rect 15596 8260 15652 8270
rect 15260 6750 15262 6802
rect 15314 6750 15316 6802
rect 15596 6916 15652 8204
rect 16044 8258 16100 8270
rect 16044 8206 16046 8258
rect 16098 8206 16100 8258
rect 16044 7924 16100 8206
rect 16044 7858 16100 7868
rect 16380 8034 16436 8046
rect 16380 7982 16382 8034
rect 16434 7982 16436 8034
rect 16380 7700 16436 7982
rect 16380 7634 16436 7644
rect 16604 7474 16660 10444
rect 16716 11956 16772 11966
rect 16716 9154 16772 11900
rect 16828 11508 16884 11518
rect 16828 10164 16884 11452
rect 16828 10098 16884 10108
rect 16716 9102 16718 9154
rect 16770 9102 16772 9154
rect 16716 9090 16772 9102
rect 16828 9716 16884 9726
rect 16828 7924 16884 9660
rect 16940 9604 16996 12348
rect 17164 11170 17220 11182
rect 17164 11118 17166 11170
rect 17218 11118 17220 11170
rect 17052 10724 17108 10734
rect 17052 10630 17108 10668
rect 17164 10612 17220 11118
rect 17276 11172 17332 12686
rect 17500 11508 17556 13020
rect 17612 12850 17668 12862
rect 17612 12798 17614 12850
rect 17666 12798 17668 12850
rect 17612 12402 17668 12798
rect 17612 12350 17614 12402
rect 17666 12350 17668 12402
rect 17612 12338 17668 12350
rect 17724 12850 17780 12862
rect 17724 12798 17726 12850
rect 17778 12798 17780 12850
rect 17500 11442 17556 11452
rect 17388 11396 17444 11406
rect 17388 11302 17444 11340
rect 17500 11284 17556 11294
rect 17500 11190 17556 11228
rect 17276 11106 17332 11116
rect 17612 11172 17668 11182
rect 17612 11078 17668 11116
rect 17612 10836 17668 10846
rect 17724 10836 17780 12798
rect 17836 12740 17892 14252
rect 18060 14196 18116 14366
rect 18172 14308 18228 14318
rect 18172 14214 18228 14252
rect 18060 14130 18116 14140
rect 18060 13860 18116 13870
rect 18060 13858 18228 13860
rect 18060 13806 18062 13858
rect 18114 13806 18228 13858
rect 18060 13804 18228 13806
rect 18060 13794 18116 13804
rect 17948 13746 18004 13758
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13188 18004 13694
rect 18172 13636 18228 13804
rect 18172 13570 18228 13580
rect 18060 13524 18116 13534
rect 18060 13430 18116 13468
rect 17948 13122 18004 13132
rect 17836 12738 18004 12740
rect 17836 12686 17838 12738
rect 17890 12686 18004 12738
rect 17836 12684 18004 12686
rect 17836 12674 17892 12684
rect 17836 12290 17892 12302
rect 17836 12238 17838 12290
rect 17890 12238 17892 12290
rect 17836 11172 17892 12238
rect 17948 12290 18004 12684
rect 17948 12238 17950 12290
rect 18002 12238 18004 12290
rect 17948 12226 18004 12238
rect 18172 12180 18228 12190
rect 18060 11620 18116 11630
rect 18060 11284 18116 11564
rect 18172 11506 18228 12124
rect 18172 11454 18174 11506
rect 18226 11454 18228 11506
rect 18172 11442 18228 11454
rect 18060 11228 18228 11284
rect 17836 11106 17892 11116
rect 17612 10834 17780 10836
rect 17612 10782 17614 10834
rect 17666 10782 17780 10834
rect 17612 10780 17780 10782
rect 17612 10770 17668 10780
rect 17836 10722 17892 10734
rect 17836 10670 17838 10722
rect 17890 10670 17892 10722
rect 17836 10612 17892 10670
rect 17164 10556 17892 10612
rect 17948 10610 18004 10622
rect 17948 10558 17950 10610
rect 18002 10558 18004 10610
rect 17052 10164 17108 10174
rect 17052 9828 17108 10108
rect 17164 10050 17220 10556
rect 17164 9998 17166 10050
rect 17218 9998 17220 10050
rect 17164 9986 17220 9998
rect 17948 10164 18004 10558
rect 17948 9940 18004 10108
rect 17948 9874 18004 9884
rect 18060 10388 18116 10398
rect 17724 9828 17780 9838
rect 17052 9772 17220 9828
rect 17052 9604 17108 9614
rect 16940 9602 17108 9604
rect 16940 9550 17054 9602
rect 17106 9550 17108 9602
rect 16940 9548 17108 9550
rect 17052 9538 17108 9548
rect 17164 8260 17220 9772
rect 17724 9734 17780 9772
rect 17836 9716 17892 9726
rect 17836 9622 17892 9660
rect 17836 9268 17892 9278
rect 17836 9174 17892 9212
rect 18060 9154 18116 10332
rect 18060 9102 18062 9154
rect 18114 9102 18116 9154
rect 18060 9090 18116 9102
rect 17612 9044 17668 9054
rect 17612 8950 17668 8988
rect 17052 8258 17220 8260
rect 17052 8206 17166 8258
rect 17218 8206 17220 8258
rect 17052 8204 17220 8206
rect 16940 8148 16996 8158
rect 16940 8054 16996 8092
rect 16828 7858 16884 7868
rect 16604 7422 16606 7474
rect 16658 7422 16660 7474
rect 16604 7410 16660 7422
rect 17052 7140 17108 8204
rect 17164 8194 17220 8204
rect 17612 8258 17668 8270
rect 17612 8206 17614 8258
rect 17666 8206 17668 8258
rect 17276 8034 17332 8046
rect 17276 7982 17278 8034
rect 17330 7982 17332 8034
rect 15596 6784 15652 6860
rect 16940 7084 17108 7140
rect 17164 7812 17220 7822
rect 16716 6804 16772 6814
rect 15260 6738 15316 6750
rect 15148 6690 15204 6702
rect 15148 6638 15150 6690
rect 15202 6638 15204 6690
rect 15148 6580 15204 6638
rect 15372 6690 15428 6702
rect 15372 6638 15374 6690
rect 15426 6638 15428 6690
rect 15260 6580 15316 6590
rect 15148 6524 15260 6580
rect 14812 5796 14868 5806
rect 14140 5742 14142 5794
rect 14194 5742 14196 5794
rect 14140 4676 14196 5742
rect 14476 5794 14868 5796
rect 14476 5742 14814 5794
rect 14866 5742 14868 5794
rect 14476 5740 14868 5742
rect 14252 5684 14308 5694
rect 14252 5682 14420 5684
rect 14252 5630 14254 5682
rect 14306 5630 14420 5682
rect 14252 5628 14420 5630
rect 14252 5618 14308 5628
rect 14252 5460 14308 5470
rect 14252 5234 14308 5404
rect 14252 5182 14254 5234
rect 14306 5182 14308 5234
rect 14252 5170 14308 5182
rect 14364 4900 14420 5628
rect 14364 4834 14420 4844
rect 14476 4676 14532 5740
rect 14812 5730 14868 5740
rect 14140 4610 14196 4620
rect 14252 4620 14532 4676
rect 14812 5236 14868 5246
rect 14028 3726 14030 3778
rect 14082 3726 14084 3778
rect 12796 3668 12852 3678
rect 12796 3574 12852 3612
rect 14028 3668 14084 3726
rect 14252 3778 14308 4620
rect 14812 4564 14868 5180
rect 15148 4788 15204 6524
rect 15260 6514 15316 6524
rect 15372 6356 15428 6638
rect 15372 6290 15428 6300
rect 15708 6690 15764 6702
rect 15708 6638 15710 6690
rect 15762 6638 15764 6690
rect 15708 6244 15764 6638
rect 16492 6690 16548 6702
rect 16492 6638 16494 6690
rect 16546 6638 16548 6690
rect 15708 6178 15764 6188
rect 16044 6578 16100 6590
rect 16044 6526 16046 6578
rect 16098 6526 16100 6578
rect 15820 6020 15876 6030
rect 15820 5926 15876 5964
rect 16044 5236 16100 6526
rect 16044 5170 16100 5180
rect 15148 4722 15204 4732
rect 15932 5010 15988 5022
rect 15932 4958 15934 5010
rect 15986 4958 15988 5010
rect 14252 3726 14254 3778
rect 14306 3726 14308 3778
rect 14252 3714 14308 3726
rect 14476 4508 14868 4564
rect 14476 3778 14532 4508
rect 14700 4340 14756 4350
rect 14700 4246 14756 4284
rect 14476 3726 14478 3778
rect 14530 3726 14532 3778
rect 14476 3714 14532 3726
rect 14028 3602 14084 3612
rect 14588 3668 14644 3678
rect 14588 3574 14644 3612
rect 15484 3668 15540 3678
rect 15484 3574 15540 3612
rect 10220 3330 10276 3342
rect 10220 3278 10222 3330
rect 10274 3278 10276 3330
rect 10220 3108 10276 3278
rect 10220 3042 10276 3052
rect 10556 3332 10612 3342
rect 10556 800 10612 3276
rect 11900 3332 12292 3388
rect 13244 3556 13300 3566
rect 11900 800 11956 3332
rect 13244 800 13300 3500
rect 13916 3442 13972 3454
rect 13916 3390 13918 3442
rect 13970 3390 13972 3442
rect 13916 2996 13972 3390
rect 14700 3444 14756 3454
rect 13916 2930 13972 2940
rect 14588 3332 14756 3388
rect 14588 800 14644 3332
rect 15932 2996 15988 4958
rect 16492 3668 16548 6638
rect 16716 5460 16772 6748
rect 16940 6692 16996 7084
rect 17052 6916 17108 6926
rect 17052 6822 17108 6860
rect 16940 6636 17108 6692
rect 16828 6578 16884 6590
rect 16828 6526 16830 6578
rect 16882 6526 16884 6578
rect 16828 6244 16884 6526
rect 16940 6468 16996 6478
rect 16940 6374 16996 6412
rect 16828 6178 16884 6188
rect 16940 6132 16996 6142
rect 16940 6038 16996 6076
rect 16828 6020 16884 6030
rect 16828 5684 16884 5964
rect 16828 5618 16884 5628
rect 16716 5394 16772 5404
rect 17052 5348 17108 6636
rect 17052 5282 17108 5292
rect 16828 5122 16884 5134
rect 16828 5070 16830 5122
rect 16882 5070 16884 5122
rect 16716 4788 16772 4798
rect 16716 4228 16772 4732
rect 16828 4452 16884 5070
rect 16828 4386 16884 4396
rect 16828 4228 16884 4238
rect 16716 4226 16884 4228
rect 16716 4174 16830 4226
rect 16882 4174 16884 4226
rect 16716 4172 16884 4174
rect 16828 4162 16884 4172
rect 16492 3602 16548 3612
rect 17164 3556 17220 7756
rect 17276 7364 17332 7982
rect 17388 8034 17444 8046
rect 17388 7982 17390 8034
rect 17442 7982 17444 8034
rect 17388 7700 17444 7982
rect 17612 7924 17668 8206
rect 17612 7868 17892 7924
rect 17612 7700 17668 7710
rect 17388 7698 17668 7700
rect 17388 7646 17614 7698
rect 17666 7646 17668 7698
rect 17388 7644 17668 7646
rect 17612 7634 17668 7644
rect 17724 7700 17780 7710
rect 17724 7606 17780 7644
rect 17276 7308 17668 7364
rect 17500 7140 17556 7150
rect 17276 6690 17332 6702
rect 17276 6638 17278 6690
rect 17330 6638 17332 6690
rect 17276 6356 17332 6638
rect 17276 6290 17332 6300
rect 17388 6692 17444 6702
rect 17388 5908 17444 6636
rect 17388 5842 17444 5852
rect 17500 6578 17556 7084
rect 17500 6526 17502 6578
rect 17554 6526 17556 6578
rect 17500 5012 17556 6526
rect 17612 5234 17668 7308
rect 17836 6468 17892 7868
rect 17948 7700 18004 7710
rect 17948 7606 18004 7644
rect 18172 7586 18228 11228
rect 18284 9154 18340 14476
rect 18396 14530 18452 15372
rect 18620 15426 18676 15484
rect 18620 15374 18622 15426
rect 18674 15374 18676 15426
rect 18620 15362 18676 15374
rect 18396 14478 18398 14530
rect 18450 14478 18452 14530
rect 18396 14466 18452 14478
rect 18508 15314 18564 15326
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 14196 18564 15262
rect 18732 15316 18788 15326
rect 18732 15222 18788 15260
rect 18508 14130 18564 14140
rect 18620 14980 18676 14990
rect 18620 13972 18676 14924
rect 18844 14084 18900 15596
rect 18508 13916 18676 13972
rect 18732 14028 18900 14084
rect 18956 15428 19012 15438
rect 18732 13972 18788 14028
rect 18508 12404 18564 13916
rect 18732 13858 18788 13916
rect 18732 13806 18734 13858
rect 18786 13806 18788 13858
rect 18732 13794 18788 13806
rect 18844 13860 18900 13870
rect 18844 13766 18900 13804
rect 18620 13748 18676 13758
rect 18620 12516 18676 13692
rect 18956 13300 19012 15372
rect 19068 14084 19124 15932
rect 19180 15540 19236 18284
rect 19292 17892 19348 17902
rect 19292 17332 19348 17836
rect 19628 17890 19684 18398
rect 20188 18340 20244 18350
rect 20188 18246 20244 18284
rect 19628 17838 19630 17890
rect 19682 17838 19684 17890
rect 19628 17826 19684 17838
rect 20300 17892 20356 18620
rect 20300 17826 20356 17836
rect 20636 18338 20692 18350
rect 20636 18286 20638 18338
rect 20690 18286 20692 18338
rect 19404 17444 19460 17454
rect 19404 17350 19460 17388
rect 19964 17444 20020 17482
rect 20412 17444 20468 17454
rect 19964 17378 20020 17388
rect 20300 17442 20468 17444
rect 20300 17390 20414 17442
rect 20466 17390 20468 17442
rect 20300 17388 20468 17390
rect 19292 17266 19348 17276
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19180 15474 19236 15484
rect 19292 17106 19908 17108
rect 19292 17054 19854 17106
rect 19906 17054 19908 17106
rect 19292 17052 19908 17054
rect 19180 15314 19236 15326
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 19180 15204 19236 15262
rect 19180 15138 19236 15148
rect 19292 14420 19348 17052
rect 19852 17042 19908 17052
rect 19740 16884 19796 16894
rect 19628 16882 19796 16884
rect 19628 16830 19742 16882
rect 19794 16830 19796 16882
rect 19628 16828 19796 16830
rect 19516 16212 19572 16222
rect 19404 15988 19460 15998
rect 19404 15894 19460 15932
rect 19516 15876 19572 16156
rect 19516 15782 19572 15820
rect 19628 15540 19684 16828
rect 19740 16818 19796 16828
rect 20076 16882 20132 16894
rect 20076 16830 20078 16882
rect 20130 16830 20132 16882
rect 20076 15988 20132 16830
rect 20076 15922 20132 15932
rect 20188 15986 20244 15998
rect 20188 15934 20190 15986
rect 20242 15934 20244 15986
rect 19740 15876 19796 15914
rect 19740 15810 19796 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19684 15484 19796 15540
rect 19628 15474 19684 15484
rect 19740 15426 19796 15484
rect 19740 15374 19742 15426
rect 19794 15374 19796 15426
rect 19740 15362 19796 15374
rect 19628 15314 19684 15326
rect 19628 15262 19630 15314
rect 19682 15262 19684 15314
rect 19516 15204 19572 15214
rect 19628 15204 19684 15262
rect 19572 15148 19684 15204
rect 19516 15138 19572 15148
rect 19404 14756 19460 14766
rect 19404 14662 19460 14700
rect 20188 14756 20244 15934
rect 20300 15540 20356 17388
rect 20412 17378 20468 17388
rect 20636 17444 20692 18286
rect 20636 17378 20692 17388
rect 20860 17892 20916 17902
rect 20860 17442 20916 17836
rect 20860 17390 20862 17442
rect 20914 17390 20916 17442
rect 20860 17220 20916 17390
rect 20860 17154 20916 17164
rect 20860 16770 20916 16782
rect 20860 16718 20862 16770
rect 20914 16718 20916 16770
rect 20748 16658 20804 16670
rect 20748 16606 20750 16658
rect 20802 16606 20804 16658
rect 20748 16322 20804 16606
rect 20748 16270 20750 16322
rect 20802 16270 20804 16322
rect 20748 16258 20804 16270
rect 20636 16212 20692 16222
rect 20412 16100 20468 16110
rect 20412 16006 20468 16044
rect 20636 15986 20692 16156
rect 20860 16212 20916 16718
rect 20860 16146 20916 16156
rect 20636 15934 20638 15986
rect 20690 15934 20692 15986
rect 20636 15652 20692 15934
rect 20636 15586 20692 15596
rect 20748 15876 20804 15886
rect 20300 15484 20468 15540
rect 20188 14690 20244 14700
rect 20300 15314 20356 15326
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 19516 14532 19572 14542
rect 19516 14438 19572 14476
rect 20076 14532 20132 14542
rect 20300 14532 20356 15262
rect 20412 15316 20468 15484
rect 20748 15538 20804 15820
rect 20748 15486 20750 15538
rect 20802 15486 20804 15538
rect 20748 15474 20804 15486
rect 20860 15540 20916 15550
rect 20860 15446 20916 15484
rect 20412 15250 20468 15260
rect 20524 15316 20580 15326
rect 20748 15316 20804 15326
rect 20524 15314 20692 15316
rect 20524 15262 20526 15314
rect 20578 15262 20692 15314
rect 20524 15260 20692 15262
rect 20524 15250 20580 15260
rect 20524 15092 20580 15102
rect 20132 14476 20356 14532
rect 20412 14532 20468 14542
rect 20076 14400 20132 14476
rect 19292 14354 19348 14364
rect 19068 13970 19124 14028
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 19068 13906 19124 13918
rect 19404 14308 19460 14318
rect 19180 13748 19236 13758
rect 18844 13244 19012 13300
rect 19068 13636 19124 13646
rect 18620 12460 18788 12516
rect 18508 12348 18676 12404
rect 18620 12290 18676 12348
rect 18620 12238 18622 12290
rect 18674 12238 18676 12290
rect 18508 12178 18564 12190
rect 18508 12126 18510 12178
rect 18562 12126 18564 12178
rect 18508 10836 18564 12126
rect 18620 11620 18676 12238
rect 18620 11554 18676 11564
rect 18732 11396 18788 12460
rect 18844 12402 18900 13244
rect 18956 12964 19012 12974
rect 19068 12964 19124 13580
rect 18956 12962 19124 12964
rect 18956 12910 18958 12962
rect 19010 12910 19124 12962
rect 18956 12908 19124 12910
rect 18956 12898 19012 12908
rect 19068 12740 19124 12750
rect 19180 12740 19236 13692
rect 19292 13412 19348 13422
rect 19404 13412 19460 14252
rect 19836 14140 20100 14150
rect 19516 14084 19572 14094
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13858 19572 14028
rect 20188 13970 20244 14476
rect 20300 14308 20356 14318
rect 20412 14308 20468 14476
rect 20524 14418 20580 15036
rect 20636 14532 20692 15260
rect 20636 14466 20692 14476
rect 20524 14366 20526 14418
rect 20578 14366 20580 14418
rect 20524 14354 20580 14366
rect 20356 14252 20468 14308
rect 20636 14308 20692 14318
rect 20300 14214 20356 14252
rect 20636 14214 20692 14252
rect 19516 13806 19518 13858
rect 19570 13806 19572 13858
rect 19516 13794 19572 13806
rect 19628 13914 19684 13926
rect 19628 13862 19630 13914
rect 19682 13862 19684 13914
rect 20188 13918 20190 13970
rect 20242 13918 20244 13970
rect 20188 13906 20244 13918
rect 20412 14084 20468 14094
rect 20412 13970 20468 14028
rect 20412 13918 20414 13970
rect 20466 13918 20468 13970
rect 20412 13906 20468 13918
rect 19628 13524 19684 13862
rect 20524 13860 20580 13870
rect 19628 13458 19684 13468
rect 19852 13746 19908 13758
rect 19852 13694 19854 13746
rect 19906 13694 19908 13746
rect 19348 13356 19460 13412
rect 19852 13412 19908 13694
rect 19292 12962 19348 13356
rect 19852 13346 19908 13356
rect 20524 13746 20580 13804
rect 20524 13694 20526 13746
rect 20578 13694 20580 13746
rect 19292 12910 19294 12962
rect 19346 12910 19348 12962
rect 19292 12898 19348 12910
rect 19516 13300 19572 13310
rect 19068 12738 19236 12740
rect 19068 12686 19070 12738
rect 19122 12686 19236 12738
rect 19068 12684 19236 12686
rect 19068 12674 19124 12684
rect 18844 12350 18846 12402
rect 18898 12350 18900 12402
rect 18844 12338 18900 12350
rect 19068 12516 19124 12526
rect 18732 11340 18900 11396
rect 18620 11282 18676 11294
rect 18620 11230 18622 11282
rect 18674 11230 18676 11282
rect 18620 11060 18676 11230
rect 18732 11172 18788 11182
rect 18732 11078 18788 11116
rect 18620 10994 18676 11004
rect 18508 10770 18564 10780
rect 18508 10612 18564 10622
rect 18508 10518 18564 10556
rect 18844 10164 18900 11340
rect 18508 10108 18900 10164
rect 18956 11170 19012 11182
rect 18956 11118 18958 11170
rect 19010 11118 19012 11170
rect 18508 9938 18564 10108
rect 18508 9886 18510 9938
rect 18562 9886 18564 9938
rect 18508 9874 18564 9886
rect 18620 9940 18676 9950
rect 18620 9826 18676 9884
rect 18956 9940 19012 11118
rect 18956 9874 19012 9884
rect 18620 9774 18622 9826
rect 18674 9774 18676 9826
rect 18620 9762 18676 9774
rect 18844 9826 18900 9838
rect 18844 9774 18846 9826
rect 18898 9774 18900 9826
rect 18284 9102 18286 9154
rect 18338 9102 18340 9154
rect 18284 9090 18340 9102
rect 18396 9714 18452 9726
rect 18396 9662 18398 9714
rect 18450 9662 18452 9714
rect 18396 8820 18452 9662
rect 18844 9604 18900 9774
rect 18844 9538 18900 9548
rect 18396 8754 18452 8764
rect 19068 8596 19124 12460
rect 19404 11396 19460 11406
rect 19404 11302 19460 11340
rect 19292 10164 19348 10174
rect 19180 9828 19236 9838
rect 19180 9266 19236 9772
rect 19180 9214 19182 9266
rect 19234 9214 19236 9266
rect 19180 9202 19236 9214
rect 19292 9266 19348 10108
rect 19516 9940 19572 13244
rect 20076 12964 20132 12974
rect 20076 12870 20132 12908
rect 20412 12962 20468 12974
rect 20412 12910 20414 12962
rect 20466 12910 20468 12962
rect 19740 12852 19796 12862
rect 19740 12758 19796 12796
rect 20188 12738 20244 12750
rect 20188 12686 20190 12738
rect 20242 12686 20244 12738
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20188 12292 20244 12686
rect 20300 12292 20356 12302
rect 20188 12290 20356 12292
rect 20188 12238 20302 12290
rect 20354 12238 20356 12290
rect 20188 12236 20356 12238
rect 20300 12226 20356 12236
rect 19628 12180 19684 12190
rect 19628 12086 19684 12124
rect 20412 11844 20468 12910
rect 20524 12292 20580 13694
rect 20524 12226 20580 12236
rect 20412 11778 20468 11788
rect 20748 11508 20804 15260
rect 20972 15148 21028 18956
rect 21084 18340 21140 18350
rect 21084 18246 21140 18284
rect 21308 17444 21364 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 42588 22596 42644 22606
rect 42252 22484 42308 22494
rect 25340 22372 25396 22382
rect 22316 22148 22372 22158
rect 21420 19906 21476 19918
rect 21420 19854 21422 19906
rect 21474 19854 21476 19906
rect 21420 19796 21476 19854
rect 21420 19730 21476 19740
rect 21532 19010 21588 19022
rect 21980 19012 22036 19022
rect 21532 18958 21534 19010
rect 21586 18958 21588 19010
rect 21532 17668 21588 18958
rect 21868 19010 22036 19012
rect 21868 18958 21982 19010
rect 22034 18958 22036 19010
rect 21868 18956 22036 18958
rect 21532 17602 21588 17612
rect 21644 18338 21700 18350
rect 21644 18286 21646 18338
rect 21698 18286 21700 18338
rect 21532 17444 21588 17454
rect 21308 17442 21588 17444
rect 21308 17390 21534 17442
rect 21586 17390 21588 17442
rect 21308 17388 21588 17390
rect 21532 17332 21588 17388
rect 21532 17266 21588 17276
rect 21644 16884 21700 18286
rect 21868 18116 21924 18956
rect 21980 18946 22036 18956
rect 22316 18676 22372 22092
rect 22540 20580 22596 20590
rect 22428 19684 22484 19694
rect 22428 19346 22484 19628
rect 22428 19294 22430 19346
rect 22482 19294 22484 19346
rect 22428 19282 22484 19294
rect 22428 18676 22484 18686
rect 22316 18674 22484 18676
rect 22316 18622 22430 18674
rect 22482 18622 22484 18674
rect 22316 18620 22484 18622
rect 22428 18610 22484 18620
rect 21868 18050 21924 18060
rect 21980 18338 22036 18350
rect 21980 18286 21982 18338
rect 22034 18286 22036 18338
rect 21644 16818 21700 16828
rect 21756 17444 21812 17454
rect 21756 16882 21812 17388
rect 21756 16830 21758 16882
rect 21810 16830 21812 16882
rect 21420 16770 21476 16782
rect 21420 16718 21422 16770
rect 21474 16718 21476 16770
rect 21420 16324 21476 16718
rect 21420 16258 21476 16268
rect 21532 16658 21588 16670
rect 21532 16606 21534 16658
rect 21586 16606 21588 16658
rect 21532 16098 21588 16606
rect 21532 16046 21534 16098
rect 21586 16046 21588 16098
rect 21532 16034 21588 16046
rect 21644 16212 21700 16222
rect 21308 15876 21364 15886
rect 21308 15538 21364 15820
rect 21308 15486 21310 15538
rect 21362 15486 21364 15538
rect 21308 15474 21364 15486
rect 21532 15652 21588 15662
rect 21532 15538 21588 15596
rect 21532 15486 21534 15538
rect 21586 15486 21588 15538
rect 21532 15474 21588 15486
rect 20860 15092 21028 15148
rect 21084 15316 21140 15326
rect 20860 13300 20916 15092
rect 20972 13636 21028 13646
rect 21084 13636 21140 15260
rect 20972 13634 21140 13636
rect 20972 13582 20974 13634
rect 21026 13582 21140 13634
rect 20972 13580 21140 13582
rect 20972 13570 21028 13580
rect 20860 13234 20916 13244
rect 21084 13300 21140 13580
rect 21084 13234 21140 13244
rect 21196 15090 21252 15102
rect 21196 15038 21198 15090
rect 21250 15038 21252 15090
rect 21196 12964 21252 15038
rect 21644 14756 21700 16156
rect 21756 14980 21812 16830
rect 21868 16324 21924 16334
rect 21868 16098 21924 16268
rect 21868 16046 21870 16098
rect 21922 16046 21924 16098
rect 21868 15316 21924 16046
rect 21868 15250 21924 15260
rect 21756 14914 21812 14924
rect 21644 14700 21812 14756
rect 21644 14530 21700 14542
rect 21644 14478 21646 14530
rect 21698 14478 21700 14530
rect 21196 12898 21252 12908
rect 21420 13972 21476 13982
rect 21420 13748 21476 13916
rect 21644 13970 21700 14478
rect 21644 13918 21646 13970
rect 21698 13918 21700 13970
rect 21644 13906 21700 13918
rect 21756 14084 21812 14700
rect 21980 14644 22036 18286
rect 22540 17778 22596 20524
rect 23548 19348 23604 19358
rect 22876 18452 22932 18462
rect 22876 18358 22932 18396
rect 22540 17726 22542 17778
rect 22594 17726 22596 17778
rect 22092 17444 22148 17454
rect 22092 17350 22148 17388
rect 22540 16884 22596 17726
rect 22652 18340 22708 18350
rect 22652 17108 22708 18284
rect 23548 17780 23604 19292
rect 23548 17648 23604 17724
rect 23100 17444 23156 17454
rect 24332 17444 24388 17454
rect 23100 17350 23156 17388
rect 24220 17442 24388 17444
rect 24220 17390 24334 17442
rect 24386 17390 24388 17442
rect 24220 17388 24388 17390
rect 22652 16976 22708 17052
rect 23548 17220 23604 17230
rect 23548 17106 23604 17164
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 22540 16828 22708 16884
rect 22204 16772 22260 16782
rect 22652 16772 22708 16828
rect 22204 16770 22372 16772
rect 22204 16718 22206 16770
rect 22258 16718 22372 16770
rect 22204 16716 22372 16718
rect 22204 16706 22260 16716
rect 22092 15874 22148 15886
rect 22092 15822 22094 15874
rect 22146 15822 22148 15874
rect 22092 15540 22148 15822
rect 22092 15474 22148 15484
rect 22204 15874 22260 15886
rect 22204 15822 22206 15874
rect 22258 15822 22260 15874
rect 22204 15428 22260 15822
rect 22204 15362 22260 15372
rect 22316 15316 22372 16716
rect 22652 16706 22708 16716
rect 23100 16770 23156 16782
rect 23100 16718 23102 16770
rect 23154 16718 23156 16770
rect 22764 16212 22820 16222
rect 22764 16118 22820 16156
rect 22652 15874 22708 15886
rect 22652 15822 22654 15874
rect 22706 15822 22708 15874
rect 22540 15316 22596 15326
rect 22316 15260 22540 15316
rect 22540 15222 22596 15260
rect 21980 14578 22036 14588
rect 21980 14420 22036 14430
rect 21980 14326 22036 14364
rect 22092 14306 22148 14318
rect 22092 14254 22094 14306
rect 22146 14254 22148 14306
rect 21756 13970 21812 14028
rect 21756 13918 21758 13970
rect 21810 13918 21812 13970
rect 21756 13906 21812 13918
rect 21980 14084 22036 14094
rect 21532 13748 21588 13758
rect 21420 13746 21588 13748
rect 21420 13694 21534 13746
rect 21586 13694 21588 13746
rect 21420 13692 21588 13694
rect 20860 12738 20916 12750
rect 20860 12686 20862 12738
rect 20914 12686 20916 12738
rect 20860 12292 20916 12686
rect 20860 12226 20916 12236
rect 20412 11452 21140 11508
rect 20412 11394 20468 11452
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20412 11330 20468 11342
rect 19628 11170 19684 11182
rect 19628 11118 19630 11170
rect 19682 11118 19684 11170
rect 19628 11060 19684 11118
rect 19852 11172 19908 11210
rect 19852 11106 19908 11116
rect 19964 11172 20020 11182
rect 20524 11172 20580 11182
rect 19964 11170 20244 11172
rect 19964 11118 19966 11170
rect 20018 11118 20244 11170
rect 19964 11116 20244 11118
rect 19964 11106 20020 11116
rect 19628 10836 19684 11004
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10780 19796 10836
rect 19292 9214 19294 9266
rect 19346 9214 19348 9266
rect 19292 9202 19348 9214
rect 19404 9884 19572 9940
rect 19628 9940 19684 9950
rect 19404 9044 19460 9884
rect 19516 9716 19572 9726
rect 19516 9622 19572 9660
rect 19628 9714 19684 9884
rect 19628 9662 19630 9714
rect 19682 9662 19684 9714
rect 19628 9650 19684 9662
rect 19740 9604 19796 10780
rect 19852 9716 19908 9726
rect 19852 9622 19908 9660
rect 19740 9538 19796 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19852 9044 19908 9054
rect 19404 8988 19684 9044
rect 19404 8820 19460 8830
rect 19404 8726 19460 8764
rect 19068 8530 19124 8540
rect 19292 8372 19348 8382
rect 19292 8258 19348 8316
rect 19516 8260 19572 8270
rect 19292 8206 19294 8258
rect 19346 8206 19348 8258
rect 18284 8148 18340 8158
rect 18284 8034 18340 8092
rect 18844 8148 18900 8158
rect 18844 8146 19012 8148
rect 18844 8094 18846 8146
rect 18898 8094 19012 8146
rect 18844 8092 19012 8094
rect 18844 8082 18900 8092
rect 18284 7982 18286 8034
rect 18338 7982 18340 8034
rect 18284 7700 18340 7982
rect 18284 7634 18340 7644
rect 18172 7534 18174 7586
rect 18226 7534 18228 7586
rect 18172 7522 18228 7534
rect 18732 7474 18788 7486
rect 18732 7422 18734 7474
rect 18786 7422 18788 7474
rect 18620 6690 18676 6702
rect 18620 6638 18622 6690
rect 18674 6638 18676 6690
rect 18396 6578 18452 6590
rect 18396 6526 18398 6578
rect 18450 6526 18452 6578
rect 18284 6468 18340 6478
rect 17836 6466 18340 6468
rect 17836 6414 18286 6466
rect 18338 6414 18340 6466
rect 17836 6412 18340 6414
rect 18284 6402 18340 6412
rect 18396 6468 18452 6526
rect 18396 6020 18452 6412
rect 18396 5954 18452 5964
rect 18508 6580 18564 6590
rect 17724 5908 17780 5918
rect 17724 5814 17780 5852
rect 18508 5796 18564 6524
rect 18620 6356 18676 6638
rect 18620 6290 18676 6300
rect 17612 5182 17614 5234
rect 17666 5182 17668 5234
rect 17612 5170 17668 5182
rect 18396 5794 18564 5796
rect 18396 5742 18510 5794
rect 18562 5742 18564 5794
rect 18396 5740 18564 5742
rect 17500 4946 17556 4956
rect 18060 5124 18116 5134
rect 17164 3490 17220 3500
rect 17612 4676 17668 4686
rect 17612 3556 17668 4620
rect 18060 4450 18116 5068
rect 18060 4398 18062 4450
rect 18114 4398 18116 4450
rect 18060 4386 18116 4398
rect 18284 4564 18340 4574
rect 18172 4340 18228 4350
rect 18172 4246 18228 4284
rect 17724 3780 17780 3790
rect 17724 3686 17780 3724
rect 16604 3442 16660 3454
rect 16604 3390 16606 3442
rect 16658 3390 16660 3442
rect 17612 3424 17668 3500
rect 18284 3554 18340 4508
rect 18396 4338 18452 5740
rect 18508 5730 18564 5740
rect 18396 4286 18398 4338
rect 18450 4286 18452 4338
rect 18396 4274 18452 4286
rect 18508 5572 18564 5582
rect 18508 4116 18564 5516
rect 18732 4452 18788 7422
rect 18844 6692 18900 6702
rect 18844 6598 18900 6636
rect 18956 4900 19012 8092
rect 19068 8146 19124 8158
rect 19068 8094 19070 8146
rect 19122 8094 19124 8146
rect 19068 7474 19124 8094
rect 19068 7422 19070 7474
rect 19122 7422 19124 7474
rect 19068 6578 19124 7422
rect 19292 7364 19348 8206
rect 19292 7298 19348 7308
rect 19404 8258 19572 8260
rect 19404 8206 19518 8258
rect 19570 8206 19572 8258
rect 19404 8204 19572 8206
rect 19404 7362 19460 8204
rect 19516 8194 19572 8204
rect 19628 7700 19684 8988
rect 19852 8930 19908 8988
rect 19852 8878 19854 8930
rect 19906 8878 19908 8930
rect 19852 8372 19908 8878
rect 19852 8306 19908 8316
rect 20188 8260 20244 11116
rect 20524 10948 20580 11116
rect 20636 11172 20692 11182
rect 20636 11170 20804 11172
rect 20636 11118 20638 11170
rect 20690 11118 20804 11170
rect 20636 11116 20804 11118
rect 20636 11106 20692 11116
rect 20524 10892 20692 10948
rect 20524 10500 20580 10510
rect 20524 10406 20580 10444
rect 20636 9826 20692 10892
rect 20636 9774 20638 9826
rect 20690 9774 20692 9826
rect 20636 9762 20692 9774
rect 20300 9714 20356 9726
rect 20300 9662 20302 9714
rect 20354 9662 20356 9714
rect 20300 9604 20356 9662
rect 20300 9538 20356 9548
rect 20412 9716 20468 9726
rect 20412 9266 20468 9660
rect 20524 9604 20580 9614
rect 20524 9510 20580 9548
rect 20412 9214 20414 9266
rect 20466 9214 20468 9266
rect 20412 8596 20468 9214
rect 20636 9268 20692 9278
rect 20636 9174 20692 9212
rect 20748 8930 20804 11116
rect 20860 11170 20916 11182
rect 20860 11118 20862 11170
rect 20914 11118 20916 11170
rect 20860 10052 20916 11118
rect 20860 9986 20916 9996
rect 20972 11170 21028 11182
rect 20972 11118 20974 11170
rect 21026 11118 21028 11170
rect 20860 9828 20916 9838
rect 20860 9734 20916 9772
rect 20748 8878 20750 8930
rect 20802 8878 20804 8930
rect 20748 8866 20804 8878
rect 20860 9042 20916 9054
rect 20860 8990 20862 9042
rect 20914 8990 20916 9042
rect 20860 8932 20916 8990
rect 20860 8866 20916 8876
rect 20412 8540 20916 8596
rect 20524 8372 20580 8382
rect 20412 8370 20580 8372
rect 20412 8318 20526 8370
rect 20578 8318 20580 8370
rect 20412 8316 20580 8318
rect 20300 8260 20356 8270
rect 20188 8258 20356 8260
rect 20188 8206 20302 8258
rect 20354 8206 20356 8258
rect 20188 8204 20356 8206
rect 20300 8194 20356 8204
rect 19740 8146 19796 8158
rect 19740 8094 19742 8146
rect 19794 8094 19796 8146
rect 19740 8036 19796 8094
rect 19740 7970 19796 7980
rect 19852 8148 19908 8158
rect 19852 8034 19908 8092
rect 19852 7982 19854 8034
rect 19906 7982 19908 8034
rect 19852 7970 19908 7982
rect 20300 8036 20356 8046
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19628 7644 19796 7700
rect 19628 7476 19684 7486
rect 19628 7382 19684 7420
rect 19404 7310 19406 7362
rect 19458 7310 19460 7362
rect 19180 7250 19236 7262
rect 19180 7198 19182 7250
rect 19234 7198 19236 7250
rect 19180 6916 19236 7198
rect 19180 6850 19236 6860
rect 19068 6526 19070 6578
rect 19122 6526 19124 6578
rect 19068 6244 19124 6526
rect 19292 6580 19348 6590
rect 19292 6486 19348 6524
rect 19404 6356 19460 7310
rect 19516 7364 19572 7374
rect 19516 7270 19572 7308
rect 19740 7252 19796 7644
rect 20300 7698 20356 7980
rect 20300 7646 20302 7698
rect 20354 7646 20356 7698
rect 20300 7634 20356 7646
rect 19404 6290 19460 6300
rect 19628 7196 19796 7252
rect 19852 7476 19908 7486
rect 19068 6178 19124 6188
rect 19628 6018 19684 7196
rect 19852 7028 19908 7420
rect 19852 6962 19908 6972
rect 20188 7364 20244 7374
rect 20188 6690 20244 7308
rect 20188 6638 20190 6690
rect 20242 6638 20244 6690
rect 20188 6626 20244 6638
rect 20412 6690 20468 8316
rect 20524 8306 20580 8316
rect 20860 8146 20916 8540
rect 20972 8484 21028 11118
rect 20972 8418 21028 8428
rect 21084 9156 21140 11452
rect 21420 11172 21476 13692
rect 21532 13682 21588 13692
rect 21980 12964 22036 14028
rect 22092 13972 22148 14254
rect 22204 14308 22260 14318
rect 22204 14214 22260 14252
rect 22092 13906 22148 13916
rect 22652 13860 22708 15822
rect 22764 15428 22820 15438
rect 22764 15334 22820 15372
rect 22988 15202 23044 15214
rect 22988 15150 22990 15202
rect 23042 15150 23044 15202
rect 22652 13794 22708 13804
rect 22764 14980 22820 14990
rect 22204 13746 22260 13758
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 13524 22260 13694
rect 22652 13636 22708 13646
rect 22652 13542 22708 13580
rect 22764 13634 22820 14924
rect 22988 14756 23044 15150
rect 22988 14690 23044 14700
rect 22764 13582 22766 13634
rect 22818 13582 22820 13634
rect 21980 12908 22148 12964
rect 21868 12852 21924 12862
rect 21868 12850 22036 12852
rect 21868 12798 21870 12850
rect 21922 12798 22036 12850
rect 21868 12796 22036 12798
rect 21868 12786 21924 12796
rect 21420 11106 21476 11116
rect 21532 12738 21588 12750
rect 21532 12686 21534 12738
rect 21586 12686 21588 12738
rect 21532 11396 21588 12686
rect 21756 12738 21812 12750
rect 21756 12686 21758 12738
rect 21810 12686 21812 12738
rect 20860 8094 20862 8146
rect 20914 8094 20916 8146
rect 20860 8082 20916 8094
rect 20636 8034 20692 8046
rect 20636 7982 20638 8034
rect 20690 7982 20692 8034
rect 20636 7924 20692 7982
rect 21084 7924 21140 9100
rect 20636 7868 21140 7924
rect 21196 11060 21252 11070
rect 21196 7812 21252 11004
rect 21420 9940 21476 9950
rect 21420 9268 21476 9884
rect 21532 9828 21588 11340
rect 21532 9762 21588 9772
rect 21644 12292 21700 12302
rect 21644 11394 21700 12236
rect 21756 11956 21812 12686
rect 21756 11890 21812 11900
rect 21980 12628 22036 12796
rect 21868 11844 21924 11854
rect 21868 11506 21924 11788
rect 21868 11454 21870 11506
rect 21922 11454 21924 11506
rect 21868 11442 21924 11454
rect 21644 11342 21646 11394
rect 21698 11342 21700 11394
rect 21420 9202 21476 9212
rect 21420 9044 21476 9054
rect 21420 8950 21476 8988
rect 20748 7756 21252 7812
rect 21420 8260 21476 8270
rect 20748 7700 20804 7756
rect 20524 7364 20580 7374
rect 20524 6802 20580 7308
rect 20524 6750 20526 6802
rect 20578 6750 20580 6802
rect 20524 6738 20580 6750
rect 20412 6638 20414 6690
rect 20466 6638 20468 6690
rect 20412 6626 20468 6638
rect 20748 6690 20804 7644
rect 20860 7476 20916 7486
rect 20860 7382 20916 7420
rect 20748 6638 20750 6690
rect 20802 6638 20804 6690
rect 20748 6626 20804 6638
rect 20636 6468 20692 6478
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20636 6132 20692 6412
rect 20636 6066 20692 6076
rect 19628 5966 19630 6018
rect 19682 5966 19684 6018
rect 18956 4844 19348 4900
rect 18732 4396 19236 4452
rect 18620 4340 18676 4350
rect 18732 4340 18788 4396
rect 18620 4338 18788 4340
rect 18620 4286 18622 4338
rect 18674 4286 18788 4338
rect 18620 4284 18788 4286
rect 18620 4274 18676 4284
rect 18508 4060 18676 4116
rect 18284 3502 18286 3554
rect 18338 3502 18340 3554
rect 18284 3490 18340 3502
rect 18508 3556 18564 3566
rect 16604 3388 16660 3390
rect 16604 3332 16884 3388
rect 15932 800 15988 2940
rect 16828 2884 16884 3332
rect 17724 3330 17780 3342
rect 17724 3278 17726 3330
rect 17778 3278 17780 3330
rect 17724 3220 17780 3278
rect 18508 3330 18564 3500
rect 18620 3554 18676 4060
rect 18732 4114 18788 4126
rect 18732 4062 18734 4114
rect 18786 4062 18788 4114
rect 18732 4004 18788 4062
rect 18732 3938 18788 3948
rect 19180 3666 19236 4396
rect 19292 4004 19348 4844
rect 19292 3938 19348 3948
rect 19516 4226 19572 4238
rect 19516 4174 19518 4226
rect 19570 4174 19572 4226
rect 19180 3614 19182 3666
rect 19234 3614 19236 3666
rect 19180 3602 19236 3614
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 3490 18676 3502
rect 19516 3556 19572 4174
rect 19516 3490 19572 3500
rect 19628 3388 19684 5966
rect 20300 5794 20356 5806
rect 20300 5742 20302 5794
rect 20354 5742 20356 5794
rect 20300 5684 20356 5742
rect 20300 5618 20356 5628
rect 20300 5348 20356 5358
rect 20300 5254 20356 5292
rect 19740 5234 19796 5246
rect 19740 5182 19742 5234
rect 19794 5182 19796 5234
rect 19740 5124 19796 5182
rect 19740 5058 19796 5068
rect 20524 5124 20580 5134
rect 20524 5030 20580 5068
rect 20188 5012 20244 5022
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18508 3278 18510 3330
rect 18562 3278 18564 3330
rect 18508 3266 18564 3278
rect 19292 3332 19684 3388
rect 20188 3442 20244 4956
rect 21420 4116 21476 8204
rect 21644 8036 21700 11342
rect 21868 11170 21924 11182
rect 21868 11118 21870 11170
rect 21922 11118 21924 11170
rect 21868 11060 21924 11118
rect 21868 10994 21924 11004
rect 21868 10052 21924 10062
rect 21868 9938 21924 9996
rect 21868 9886 21870 9938
rect 21922 9886 21924 9938
rect 21868 9874 21924 9886
rect 21980 9940 22036 12572
rect 22092 11170 22148 12908
rect 22204 12292 22260 13468
rect 22764 13524 22820 13582
rect 22764 13458 22820 13468
rect 22988 14530 23044 14542
rect 22988 14478 22990 14530
rect 23042 14478 23044 14530
rect 22652 13412 22708 13422
rect 22540 13188 22596 13198
rect 22540 12850 22596 13132
rect 22540 12798 22542 12850
rect 22594 12798 22596 12850
rect 22540 12786 22596 12798
rect 22652 12850 22708 13356
rect 22876 13300 22932 13310
rect 22652 12798 22654 12850
rect 22706 12798 22708 12850
rect 22316 12740 22372 12750
rect 22316 12646 22372 12684
rect 22540 12516 22596 12526
rect 22316 12292 22372 12302
rect 22204 12236 22316 12292
rect 22316 12068 22372 12236
rect 22428 12068 22484 12078
rect 22316 12066 22484 12068
rect 22316 12014 22430 12066
rect 22482 12014 22484 12066
rect 22316 12012 22484 12014
rect 22428 12002 22484 12012
rect 22092 11118 22094 11170
rect 22146 11118 22148 11170
rect 22092 10724 22148 11118
rect 22092 10658 22148 10668
rect 22204 11396 22260 11406
rect 22204 10612 22260 11340
rect 22540 10836 22596 12460
rect 22652 11844 22708 12798
rect 22652 11778 22708 11788
rect 22764 12964 22820 12974
rect 22764 11396 22820 12908
rect 22204 10546 22260 10556
rect 22316 10780 22596 10836
rect 22652 11340 22820 11396
rect 21980 9874 22036 9884
rect 21644 7970 21700 7980
rect 21756 9602 21812 9614
rect 21756 9550 21758 9602
rect 21810 9550 21812 9602
rect 21532 7364 21588 7374
rect 21532 7270 21588 7308
rect 21756 6804 21812 9550
rect 21980 9604 22036 9614
rect 21980 9510 22036 9548
rect 22092 9042 22148 9054
rect 22092 8990 22094 9042
rect 22146 8990 22148 9042
rect 21980 8596 22036 8606
rect 21980 8370 22036 8540
rect 21980 8318 21982 8370
rect 22034 8318 22036 8370
rect 21980 8306 22036 8318
rect 21868 8148 21924 8158
rect 21868 8054 21924 8092
rect 21756 6738 21812 6748
rect 22092 7476 22148 8990
rect 22204 8484 22260 8494
rect 22204 8258 22260 8428
rect 22204 8206 22206 8258
rect 22258 8206 22260 8258
rect 22204 8194 22260 8206
rect 21868 6692 21924 6702
rect 22092 6692 22148 7420
rect 22092 6636 22260 6692
rect 21644 6466 21700 6478
rect 21644 6414 21646 6466
rect 21698 6414 21700 6466
rect 21644 6356 21700 6414
rect 21644 5460 21700 6300
rect 21756 6466 21812 6478
rect 21756 6414 21758 6466
rect 21810 6414 21812 6466
rect 21756 6020 21812 6414
rect 21756 5954 21812 5964
rect 21868 6466 21924 6636
rect 21868 6414 21870 6466
rect 21922 6414 21924 6466
rect 21868 5908 21924 6414
rect 21868 5842 21924 5852
rect 21644 5124 21700 5404
rect 22204 5124 22260 6636
rect 22316 6690 22372 10780
rect 22652 10052 22708 11340
rect 22764 11172 22820 11182
rect 22764 10388 22820 11116
rect 22764 10322 22820 10332
rect 22652 9986 22708 9996
rect 22876 9938 22932 13244
rect 22876 9886 22878 9938
rect 22930 9886 22932 9938
rect 22876 9874 22932 9886
rect 22988 12180 23044 14478
rect 23100 12964 23156 16718
rect 23212 16212 23268 16222
rect 23212 15876 23268 16156
rect 23996 15876 24052 15886
rect 23212 15810 23268 15820
rect 23884 15874 24052 15876
rect 23884 15822 23998 15874
rect 24050 15822 24052 15874
rect 23884 15820 24052 15822
rect 23884 15428 23940 15820
rect 23996 15810 24052 15820
rect 23212 15316 23268 15326
rect 23212 15222 23268 15260
rect 23772 15202 23828 15214
rect 23772 15150 23774 15202
rect 23826 15150 23828 15202
rect 23660 15090 23716 15102
rect 23660 15038 23662 15090
rect 23714 15038 23716 15090
rect 23660 14084 23716 15038
rect 23772 14980 23828 15150
rect 23884 15148 23940 15372
rect 24220 15148 24276 17388
rect 24332 17378 24388 17388
rect 23884 15092 24052 15148
rect 23772 14914 23828 14924
rect 23996 14868 24052 15092
rect 23772 14756 23828 14766
rect 23772 14642 23828 14700
rect 23772 14590 23774 14642
rect 23826 14590 23828 14642
rect 23772 14578 23828 14590
rect 23660 14028 23940 14084
rect 23324 13972 23380 13982
rect 23324 13858 23380 13916
rect 23884 13860 23940 14028
rect 23324 13806 23326 13858
rect 23378 13806 23380 13858
rect 23324 13794 23380 13806
rect 23548 13804 23884 13860
rect 23548 13746 23604 13804
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 23884 13728 23940 13804
rect 23548 13682 23604 13694
rect 23100 12898 23156 12908
rect 23324 13524 23380 13534
rect 23324 12962 23380 13468
rect 23884 13522 23940 13534
rect 23884 13470 23886 13522
rect 23938 13470 23940 13522
rect 23324 12910 23326 12962
rect 23378 12910 23380 12962
rect 23324 12898 23380 12910
rect 23548 13300 23604 13310
rect 23548 12962 23604 13244
rect 23884 13076 23940 13470
rect 23548 12910 23550 12962
rect 23602 12910 23604 12962
rect 23548 12898 23604 12910
rect 23772 13020 23940 13076
rect 23772 12850 23828 13020
rect 23772 12798 23774 12850
rect 23826 12798 23828 12850
rect 23772 12786 23828 12798
rect 23100 12740 23156 12750
rect 23100 12290 23156 12684
rect 23884 12738 23940 12750
rect 23884 12686 23886 12738
rect 23938 12686 23940 12738
rect 23772 12516 23828 12526
rect 23212 12404 23268 12442
rect 23212 12338 23268 12348
rect 23492 12404 23548 12424
rect 23548 12348 23604 12404
rect 23492 12338 23604 12348
rect 23100 12238 23102 12290
rect 23154 12238 23156 12290
rect 23100 12226 23156 12238
rect 22428 9826 22484 9838
rect 22428 9774 22430 9826
rect 22482 9774 22484 9826
rect 22428 8372 22484 9774
rect 22988 9828 23044 12124
rect 23324 12178 23380 12190
rect 23324 12126 23326 12178
rect 23378 12126 23380 12178
rect 23100 12068 23156 12078
rect 23324 12068 23380 12126
rect 23436 12180 23492 12190
rect 23436 12086 23492 12124
rect 23156 12012 23268 12068
rect 23100 12002 23156 12012
rect 22988 9762 23044 9772
rect 23100 10500 23156 10510
rect 22764 8930 22820 8942
rect 22764 8878 22766 8930
rect 22818 8878 22820 8930
rect 22764 8596 22820 8878
rect 22764 8530 22820 8540
rect 22428 8306 22484 8316
rect 23100 8258 23156 10444
rect 23100 8206 23102 8258
rect 23154 8206 23156 8258
rect 22428 8146 22484 8158
rect 22428 8094 22430 8146
rect 22482 8094 22484 8146
rect 22428 7700 22484 8094
rect 22428 7634 22484 7644
rect 23100 6916 23156 8206
rect 23100 6850 23156 6860
rect 22316 6638 22318 6690
rect 22370 6638 22372 6690
rect 22316 6626 22372 6638
rect 23212 6132 23268 12012
rect 23324 12002 23380 12012
rect 23548 11732 23604 12338
rect 23548 11394 23604 11676
rect 23660 12292 23716 12302
rect 23660 11620 23716 12236
rect 23660 11554 23716 11564
rect 23772 11396 23828 12460
rect 23884 11956 23940 12686
rect 23996 12516 24052 14812
rect 23996 12450 24052 12460
rect 24108 15092 24276 15148
rect 24332 17108 24388 17118
rect 24108 12180 24164 15092
rect 24332 13412 24388 17052
rect 24780 16996 24836 17006
rect 24780 16902 24836 16940
rect 24892 15874 24948 15886
rect 24892 15822 24894 15874
rect 24946 15822 24948 15874
rect 24556 15540 24612 15550
rect 24444 15428 24500 15438
rect 24444 15334 24500 15372
rect 24556 15426 24612 15484
rect 24892 15540 24948 15822
rect 25228 15876 25284 15886
rect 25228 15782 25284 15820
rect 24892 15474 24948 15484
rect 24556 15374 24558 15426
rect 24610 15374 24612 15426
rect 24556 15362 24612 15374
rect 24668 15428 24724 15438
rect 24668 15148 24724 15372
rect 25228 15316 25284 15326
rect 24444 15092 24836 15148
rect 24444 15090 24500 15092
rect 24444 15038 24446 15090
rect 24498 15038 24500 15090
rect 24444 15026 24500 15038
rect 24556 13972 24612 13982
rect 24556 13878 24612 13916
rect 24444 13860 24500 13870
rect 24444 13766 24500 13804
rect 24556 13524 24612 13534
rect 24556 13430 24612 13468
rect 24332 13346 24388 13356
rect 24668 13412 24724 13422
rect 24220 13076 24276 13086
rect 24220 12402 24276 13020
rect 24220 12350 24222 12402
rect 24274 12350 24276 12402
rect 24220 12338 24276 12350
rect 24444 13076 24500 13086
rect 24444 12180 24500 13020
rect 24668 12964 24724 13356
rect 24556 12962 24724 12964
rect 24556 12910 24670 12962
rect 24722 12910 24724 12962
rect 24556 12908 24724 12910
rect 24556 12740 24612 12908
rect 24668 12898 24724 12908
rect 24780 12740 24836 15092
rect 24556 12674 24612 12684
rect 24668 12684 24836 12740
rect 25004 12738 25060 12750
rect 25004 12686 25006 12738
rect 25058 12686 25060 12738
rect 24556 12180 24612 12190
rect 24444 12178 24612 12180
rect 24444 12126 24558 12178
rect 24610 12126 24612 12178
rect 24444 12124 24612 12126
rect 24108 12114 24164 12124
rect 24444 11956 24500 11966
rect 23884 11900 24388 11956
rect 23548 11342 23550 11394
rect 23602 11342 23604 11394
rect 23548 11330 23604 11342
rect 23660 11340 23828 11396
rect 23884 11620 23940 11630
rect 23884 11394 23940 11564
rect 23884 11342 23886 11394
rect 23938 11342 23940 11394
rect 23660 11170 23716 11340
rect 23884 11330 23940 11342
rect 23996 11396 24052 11406
rect 23996 11302 24052 11340
rect 23660 11118 23662 11170
rect 23714 11118 23716 11170
rect 23436 9828 23492 9838
rect 23548 9828 23604 9838
rect 23436 9826 23548 9828
rect 23436 9774 23438 9826
rect 23490 9774 23548 9826
rect 23436 9772 23548 9774
rect 23436 9762 23492 9772
rect 23436 9268 23492 9278
rect 23212 6076 23380 6132
rect 22428 6020 22484 6030
rect 22428 5926 22484 5964
rect 22988 5908 23044 5918
rect 21644 5068 21812 5124
rect 21756 5012 21812 5068
rect 22204 5058 22260 5068
rect 22540 5124 22596 5134
rect 21868 5012 21924 5022
rect 21756 5010 21924 5012
rect 21756 4958 21870 5010
rect 21922 4958 21924 5010
rect 21756 4956 21924 4958
rect 21644 4452 21700 4462
rect 21644 4358 21700 4396
rect 21420 4050 21476 4060
rect 21532 4004 21588 4014
rect 21532 3666 21588 3948
rect 21868 3892 21924 4956
rect 22428 5012 22484 5022
rect 22428 4918 22484 4956
rect 22092 4900 22148 4910
rect 22092 4806 22148 4844
rect 22204 4898 22260 4910
rect 22204 4846 22206 4898
rect 22258 4846 22260 4898
rect 22204 4452 22260 4846
rect 22204 4386 22260 4396
rect 22316 4898 22372 4910
rect 22316 4846 22318 4898
rect 22370 4846 22372 4898
rect 22316 4676 22372 4846
rect 21868 3826 21924 3836
rect 22316 3780 22372 4620
rect 22428 4340 22484 4350
rect 22540 4340 22596 5068
rect 22988 4564 23044 5852
rect 23212 5906 23268 5918
rect 23212 5854 23214 5906
rect 23266 5854 23268 5906
rect 23212 5124 23268 5854
rect 23212 5058 23268 5068
rect 23100 5010 23156 5022
rect 23100 4958 23102 5010
rect 23154 4958 23156 5010
rect 23100 4788 23156 4958
rect 23100 4722 23156 4732
rect 23212 4898 23268 4910
rect 23212 4846 23214 4898
rect 23266 4846 23268 4898
rect 22988 4498 23044 4508
rect 23212 4564 23268 4846
rect 23212 4498 23268 4508
rect 22428 4338 22596 4340
rect 22428 4286 22430 4338
rect 22482 4286 22596 4338
rect 22428 4284 22596 4286
rect 22428 4274 22484 4284
rect 22316 3714 22372 3724
rect 23100 4226 23156 4238
rect 23100 4174 23102 4226
rect 23154 4174 23156 4226
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 20188 3390 20190 3442
rect 20242 3390 20244 3442
rect 17724 3154 17780 3164
rect 16828 2818 16884 2828
rect 17276 2884 17332 2894
rect 17276 800 17332 2828
rect 18620 924 18900 980
rect 18620 800 18676 924
rect 1120 0 1232 800
rect 2464 0 2576 800
rect 3808 0 3920 800
rect 5152 0 5264 800
rect 6496 0 6608 800
rect 7840 0 7952 800
rect 9184 0 9296 800
rect 10528 0 10640 800
rect 11872 0 11984 800
rect 13216 0 13328 800
rect 14560 0 14672 800
rect 15904 0 16016 800
rect 17248 0 17360 800
rect 18592 0 18704 800
rect 18844 756 18900 924
rect 19292 756 19348 3332
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 2996 20244 3390
rect 19964 2940 20244 2996
rect 21308 3444 21364 3454
rect 19964 800 20020 2940
rect 21308 800 21364 3388
rect 22540 3444 22596 3482
rect 23100 3388 23156 4174
rect 22540 3378 22596 3388
rect 22652 3332 23156 3388
rect 23324 3444 23380 6076
rect 23436 5122 23492 9212
rect 23548 6802 23604 9772
rect 23660 9044 23716 11118
rect 23772 11170 23828 11182
rect 23772 11118 23774 11170
rect 23826 11118 23828 11170
rect 23772 11060 23828 11118
rect 24332 11172 24388 11900
rect 24444 11396 24500 11900
rect 24556 11732 24612 12124
rect 24556 11666 24612 11676
rect 24556 11396 24612 11406
rect 24444 11394 24612 11396
rect 24444 11342 24558 11394
rect 24610 11342 24612 11394
rect 24444 11340 24612 11342
rect 24556 11330 24612 11340
rect 24332 11116 24612 11172
rect 23772 11004 24276 11060
rect 23884 10836 23940 10846
rect 23660 8978 23716 8988
rect 23772 10052 23828 10062
rect 23660 7364 23716 7374
rect 23660 7270 23716 7308
rect 23548 6750 23550 6802
rect 23602 6750 23604 6802
rect 23548 6738 23604 6750
rect 23772 6130 23828 9996
rect 23772 6078 23774 6130
rect 23826 6078 23828 6130
rect 23772 6066 23828 6078
rect 23884 8148 23940 10780
rect 24220 10610 24276 11004
rect 24220 10558 24222 10610
rect 24274 10558 24276 10610
rect 24220 10546 24276 10558
rect 24556 10610 24612 11116
rect 24556 10558 24558 10610
rect 24610 10558 24612 10610
rect 24556 10546 24612 10558
rect 24444 10498 24500 10510
rect 24444 10446 24446 10498
rect 24498 10446 24500 10498
rect 24444 10164 24500 10446
rect 24108 10108 24500 10164
rect 24556 10388 24612 10398
rect 24108 9938 24164 10108
rect 24108 9886 24110 9938
rect 24162 9886 24164 9938
rect 24108 9874 24164 9886
rect 24556 8820 24612 10332
rect 23884 5908 23940 8092
rect 24220 8596 24276 8606
rect 24220 7474 24276 8540
rect 24444 7700 24500 7710
rect 24444 7606 24500 7644
rect 24220 7422 24222 7474
rect 24274 7422 24276 7474
rect 24220 6692 24276 7422
rect 24556 7250 24612 8764
rect 24556 7198 24558 7250
rect 24610 7198 24612 7250
rect 24556 7028 24612 7198
rect 24556 6962 24612 6972
rect 24220 6626 24276 6636
rect 24332 6916 24388 6926
rect 23436 5070 23438 5122
rect 23490 5070 23492 5122
rect 23436 5058 23492 5070
rect 23772 5852 23940 5908
rect 24220 6356 24276 6366
rect 24220 5908 24276 6300
rect 23548 3892 23604 3902
rect 23548 3778 23604 3836
rect 23548 3726 23550 3778
rect 23602 3726 23604 3778
rect 23548 3714 23604 3726
rect 23324 3378 23380 3388
rect 23772 3442 23828 5852
rect 24220 5814 24276 5852
rect 23996 5124 24052 5134
rect 23996 5030 24052 5068
rect 23996 4338 24052 4350
rect 23996 4286 23998 4338
rect 24050 4286 24052 4338
rect 23884 3780 23940 3790
rect 23996 3780 24052 4286
rect 23884 3778 24052 3780
rect 23884 3726 23886 3778
rect 23938 3726 24052 3778
rect 23884 3724 24052 3726
rect 23884 3714 23940 3724
rect 24332 3668 24388 6860
rect 24444 6132 24500 6142
rect 24668 6132 24724 12684
rect 25004 12404 25060 12686
rect 25004 12338 25060 12348
rect 24780 12068 24836 12078
rect 24780 12066 25172 12068
rect 24780 12014 24782 12066
rect 24834 12014 25172 12066
rect 24780 12012 25172 12014
rect 24780 12002 24836 12012
rect 24892 11844 24948 11854
rect 24892 11508 24948 11788
rect 25116 11620 25172 12012
rect 25116 11554 25172 11564
rect 24780 11452 24948 11508
rect 24780 11170 24836 11452
rect 25004 11396 25060 11406
rect 24892 11284 24948 11294
rect 24892 11190 24948 11228
rect 24780 11118 24782 11170
rect 24834 11118 24836 11170
rect 24780 6468 24836 11118
rect 24892 10610 24948 10622
rect 24892 10558 24894 10610
rect 24946 10558 24948 10610
rect 24892 10052 24948 10558
rect 25004 10276 25060 11340
rect 25004 10210 25060 10220
rect 24892 9986 24948 9996
rect 24892 8930 24948 8942
rect 24892 8878 24894 8930
rect 24946 8878 24948 8930
rect 24892 8820 24948 8878
rect 25228 8932 25284 15260
rect 25340 15148 25396 22316
rect 39116 22372 39172 22382
rect 39116 22278 39172 22316
rect 40572 22372 40628 22382
rect 40012 22258 40068 22270
rect 40012 22206 40014 22258
rect 40066 22206 40068 22258
rect 40012 22036 40068 22206
rect 40012 21970 40068 21980
rect 40572 22146 40628 22316
rect 40572 22094 40574 22146
rect 40626 22094 40628 22146
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 26908 17442 26964 17454
rect 26908 17390 26910 17442
rect 26962 17390 26964 17442
rect 26460 16884 26516 16894
rect 26460 16790 26516 16828
rect 25676 16772 25732 16782
rect 25676 16770 25956 16772
rect 25676 16718 25678 16770
rect 25730 16718 25956 16770
rect 25676 16716 25956 16718
rect 25676 16706 25732 16716
rect 25676 15428 25732 15438
rect 25676 15334 25732 15372
rect 25788 15204 25844 15242
rect 25340 15092 25620 15148
rect 25788 15138 25844 15148
rect 25452 14980 25508 14990
rect 25340 14868 25396 14878
rect 25340 11508 25396 14812
rect 25452 12404 25508 14924
rect 25564 13860 25620 15092
rect 25900 14868 25956 16716
rect 26124 16770 26180 16782
rect 26124 16718 26126 16770
rect 26178 16718 26180 16770
rect 26012 15874 26068 15886
rect 26012 15822 26014 15874
rect 26066 15822 26068 15874
rect 26012 15092 26068 15822
rect 26124 15540 26180 16718
rect 26460 15874 26516 15886
rect 26796 15876 26852 15886
rect 26460 15822 26462 15874
rect 26514 15822 26516 15874
rect 26236 15540 26292 15550
rect 26124 15538 26292 15540
rect 26124 15486 26238 15538
rect 26290 15486 26292 15538
rect 26124 15484 26292 15486
rect 26124 15428 26180 15484
rect 26236 15474 26292 15484
rect 26124 15362 26180 15372
rect 26460 15148 26516 15822
rect 26684 15874 26852 15876
rect 26684 15822 26798 15874
rect 26850 15822 26852 15874
rect 26684 15820 26852 15822
rect 26684 15316 26740 15820
rect 26796 15810 26852 15820
rect 26684 15250 26740 15260
rect 26012 15026 26068 15036
rect 26124 15092 26516 15148
rect 26796 15202 26852 15214
rect 26796 15150 26798 15202
rect 26850 15150 26852 15202
rect 25900 14812 26068 14868
rect 25900 14644 25956 14654
rect 25564 13794 25620 13804
rect 25788 14642 25956 14644
rect 25788 14590 25902 14642
rect 25954 14590 25956 14642
rect 25788 14588 25956 14590
rect 25564 13636 25620 13646
rect 25788 13636 25844 14588
rect 25900 14578 25956 14588
rect 26012 14420 26068 14812
rect 26012 14354 26068 14364
rect 26012 13748 26068 13758
rect 25564 13634 25844 13636
rect 25564 13582 25566 13634
rect 25618 13582 25844 13634
rect 25564 13580 25844 13582
rect 25900 13692 26012 13748
rect 25564 13412 25620 13580
rect 25564 13346 25620 13356
rect 25564 13188 25620 13198
rect 25564 13094 25620 13132
rect 25676 12850 25732 12862
rect 25676 12798 25678 12850
rect 25730 12798 25732 12850
rect 25676 12628 25732 12798
rect 25676 12562 25732 12572
rect 25564 12404 25620 12414
rect 25452 12402 25620 12404
rect 25452 12350 25566 12402
rect 25618 12350 25620 12402
rect 25452 12348 25620 12350
rect 25564 12338 25620 12348
rect 25788 12404 25844 12414
rect 25788 12310 25844 12348
rect 25900 12290 25956 13692
rect 26012 13616 26068 13692
rect 25900 12238 25902 12290
rect 25954 12238 25956 12290
rect 25900 12226 25956 12238
rect 25340 11442 25396 11452
rect 25676 11732 25732 11742
rect 25676 11394 25732 11676
rect 25676 11342 25678 11394
rect 25730 11342 25732 11394
rect 25676 10164 25732 11342
rect 25788 11620 25844 11630
rect 25788 11282 25844 11564
rect 26012 11396 26068 11406
rect 26012 11302 26068 11340
rect 25788 11230 25790 11282
rect 25842 11230 25844 11282
rect 25788 11218 25844 11230
rect 25900 11172 25956 11182
rect 25676 10098 25732 10108
rect 25788 10388 25844 10398
rect 25228 8866 25284 8876
rect 25676 8930 25732 8942
rect 25676 8878 25678 8930
rect 25730 8878 25732 8930
rect 24892 8754 24948 8764
rect 24780 6402 24836 6412
rect 24892 8484 24948 8494
rect 24780 6132 24836 6142
rect 24668 6130 24836 6132
rect 24668 6078 24782 6130
rect 24834 6078 24836 6130
rect 24668 6076 24836 6078
rect 24444 6038 24500 6076
rect 24780 6066 24836 6076
rect 24668 5908 24724 5918
rect 24892 5908 24948 8428
rect 24668 5906 24948 5908
rect 24668 5854 24670 5906
rect 24722 5854 24948 5906
rect 24668 5852 24948 5854
rect 25564 7924 25620 7934
rect 25564 6804 25620 7868
rect 25676 7588 25732 8878
rect 25788 7698 25844 10332
rect 25900 8820 25956 11116
rect 26124 11172 26180 15092
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 13972 26404 14254
rect 26348 13906 26404 13916
rect 26460 14306 26516 14318
rect 26460 14254 26462 14306
rect 26514 14254 26516 14306
rect 26348 13748 26404 13758
rect 26460 13748 26516 14254
rect 26684 14308 26740 14318
rect 26684 14214 26740 14252
rect 26348 13746 26516 13748
rect 26348 13694 26350 13746
rect 26402 13694 26516 13746
rect 26348 13692 26516 13694
rect 26572 13860 26628 13870
rect 26236 13634 26292 13646
rect 26236 13582 26238 13634
rect 26290 13582 26292 13634
rect 26236 12962 26292 13582
rect 26348 13524 26404 13692
rect 26348 13458 26404 13468
rect 26236 12910 26238 12962
rect 26290 12910 26292 12962
rect 26236 12898 26292 12910
rect 26460 12964 26516 12974
rect 26460 12870 26516 12908
rect 26348 12738 26404 12750
rect 26348 12686 26350 12738
rect 26402 12686 26404 12738
rect 26348 12516 26404 12686
rect 26348 12450 26404 12460
rect 26572 12292 26628 13804
rect 26684 13746 26740 13758
rect 26684 13694 26686 13746
rect 26738 13694 26740 13746
rect 26684 13524 26740 13694
rect 26684 13458 26740 13468
rect 26796 13636 26852 15150
rect 26908 15204 26964 17390
rect 27804 16996 27860 17006
rect 27356 16994 27860 16996
rect 27356 16942 27806 16994
rect 27858 16942 27860 16994
rect 27356 16940 27860 16942
rect 27020 16770 27076 16782
rect 27020 16718 27022 16770
rect 27074 16718 27076 16770
rect 27020 16658 27076 16718
rect 27020 16606 27022 16658
rect 27074 16606 27076 16658
rect 27020 16594 27076 16606
rect 26908 15138 26964 15148
rect 27132 15876 27188 15886
rect 27132 15538 27188 15820
rect 27132 15486 27134 15538
rect 27186 15486 27188 15538
rect 27132 15148 27188 15486
rect 27244 15874 27300 15886
rect 27244 15822 27246 15874
rect 27298 15822 27300 15874
rect 27244 15316 27300 15822
rect 27244 15250 27300 15260
rect 27132 15092 27300 15148
rect 26124 11106 26180 11116
rect 26348 12236 26628 12292
rect 26348 11170 26404 12236
rect 26684 12180 26740 12190
rect 26796 12180 26852 13580
rect 27020 14530 27076 14542
rect 27020 14478 27022 14530
rect 27074 14478 27076 14530
rect 27020 13524 27076 14478
rect 27132 14308 27188 14318
rect 27132 13748 27188 14252
rect 27244 14196 27300 15092
rect 27356 14308 27412 16940
rect 27804 16930 27860 16940
rect 27468 16772 27524 16782
rect 27468 16678 27524 16716
rect 29484 16772 29540 16782
rect 27692 16658 27748 16670
rect 27692 16606 27694 16658
rect 27746 16606 27748 16658
rect 27468 16548 27524 16558
rect 27468 14644 27524 16492
rect 27692 15876 27748 16606
rect 29484 16212 29540 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 29932 16212 29988 16222
rect 29484 16210 29932 16212
rect 29484 16158 29486 16210
rect 29538 16158 29932 16210
rect 29484 16156 29932 16158
rect 29484 16146 29540 16156
rect 29932 16080 29988 16156
rect 34300 16212 34356 16222
rect 27692 15874 27860 15876
rect 27692 15822 27694 15874
rect 27746 15822 27860 15874
rect 27692 15820 27860 15822
rect 27692 15810 27748 15820
rect 27580 15204 27636 15214
rect 27580 15202 27748 15204
rect 27580 15150 27582 15202
rect 27634 15150 27748 15202
rect 27580 15148 27748 15150
rect 27580 15138 27636 15148
rect 27468 14550 27524 14588
rect 27580 14308 27636 14318
rect 27356 14252 27580 14308
rect 27580 14214 27636 14252
rect 27244 14140 27524 14196
rect 27356 13860 27412 13870
rect 27132 13654 27188 13692
rect 27244 13858 27412 13860
rect 27244 13806 27358 13858
rect 27410 13806 27412 13858
rect 27244 13804 27412 13806
rect 27020 13458 27076 13468
rect 27244 13076 27300 13804
rect 27356 13794 27412 13804
rect 27468 13748 27524 14140
rect 27468 13746 27636 13748
rect 27468 13694 27470 13746
rect 27522 13694 27636 13746
rect 27468 13692 27636 13694
rect 27468 13682 27524 13692
rect 27468 13524 27524 13534
rect 27468 13186 27524 13468
rect 27468 13134 27470 13186
rect 27522 13134 27524 13186
rect 27468 13122 27524 13134
rect 27244 13010 27300 13020
rect 26684 12178 26852 12180
rect 26684 12126 26686 12178
rect 26738 12126 26852 12178
rect 26684 12124 26852 12126
rect 26908 12962 26964 12974
rect 26908 12910 26910 12962
rect 26962 12910 26964 12962
rect 26684 11732 26740 12124
rect 26908 12068 26964 12910
rect 27356 12850 27412 12862
rect 27356 12798 27358 12850
rect 27410 12798 27412 12850
rect 26908 12002 26964 12012
rect 27020 12180 27076 12190
rect 26796 11956 26852 11966
rect 26796 11788 26852 11900
rect 26796 11732 26964 11788
rect 26348 11118 26350 11170
rect 26402 11118 26404 11170
rect 26348 10948 26404 11118
rect 26124 10892 26404 10948
rect 26460 11676 26740 11732
rect 26012 10610 26068 10622
rect 26012 10558 26014 10610
rect 26066 10558 26068 10610
rect 26012 9828 26068 10558
rect 26012 9044 26068 9772
rect 26012 8978 26068 8988
rect 25900 8764 26068 8820
rect 25788 7646 25790 7698
rect 25842 7646 25844 7698
rect 25788 7634 25844 7646
rect 25676 7522 25732 7532
rect 25900 7586 25956 7598
rect 25900 7534 25902 7586
rect 25954 7534 25956 7586
rect 25788 7476 25844 7486
rect 25564 5908 25620 6748
rect 25676 7250 25732 7262
rect 25676 7198 25678 7250
rect 25730 7198 25732 7250
rect 25676 6580 25732 7198
rect 25676 6132 25732 6524
rect 25676 6066 25732 6076
rect 25676 5908 25732 5918
rect 25564 5906 25732 5908
rect 25564 5854 25678 5906
rect 25730 5854 25732 5906
rect 25564 5852 25732 5854
rect 24668 5842 24724 5852
rect 25676 5842 25732 5852
rect 24556 5794 24612 5806
rect 24556 5742 24558 5794
rect 24610 5742 24612 5794
rect 24556 5348 24612 5742
rect 24556 5282 24612 5292
rect 24780 5684 24836 5694
rect 24668 5236 24724 5246
rect 24668 5142 24724 5180
rect 24780 4450 24836 5628
rect 24780 4398 24782 4450
rect 24834 4398 24836 4450
rect 24780 4386 24836 4398
rect 25788 5124 25844 7420
rect 25900 6356 25956 7534
rect 25900 6290 25956 6300
rect 25788 4338 25844 5068
rect 25788 4286 25790 4338
rect 25842 4286 25844 4338
rect 25788 4274 25844 4286
rect 24892 4114 24948 4126
rect 24892 4062 24894 4114
rect 24946 4062 24948 4114
rect 24892 3892 24948 4062
rect 24892 3826 24948 3836
rect 24444 3668 24500 3678
rect 24332 3666 24500 3668
rect 24332 3614 24446 3666
rect 24498 3614 24500 3666
rect 24332 3612 24500 3614
rect 24444 3602 24500 3612
rect 25340 3668 25396 3678
rect 23772 3390 23774 3442
rect 23826 3390 23828 3442
rect 23772 3378 23828 3390
rect 23996 3444 24052 3454
rect 22652 800 22708 3332
rect 23996 800 24052 3388
rect 25340 800 25396 3612
rect 25452 3444 25508 3482
rect 26012 3388 26068 8764
rect 26124 8260 26180 10892
rect 26236 10164 26292 10174
rect 26236 9938 26292 10108
rect 26236 9886 26238 9938
rect 26290 9886 26292 9938
rect 26236 9874 26292 9886
rect 26460 9828 26516 11676
rect 26684 11508 26740 11518
rect 26684 11394 26740 11452
rect 26684 11342 26686 11394
rect 26738 11342 26740 11394
rect 26684 11330 26740 11342
rect 26572 11172 26628 11182
rect 26572 11078 26628 11116
rect 26796 10500 26852 10510
rect 26796 10406 26852 10444
rect 26684 10276 26740 10286
rect 26684 9938 26740 10220
rect 26684 9886 26686 9938
rect 26738 9886 26740 9938
rect 26684 9874 26740 9886
rect 26460 9762 26516 9772
rect 26348 9492 26404 9502
rect 26124 8194 26180 8204
rect 26236 8932 26292 8942
rect 26236 7364 26292 8876
rect 26236 7298 26292 7308
rect 26236 6692 26292 6702
rect 26236 5906 26292 6636
rect 26236 5854 26238 5906
rect 26290 5854 26292 5906
rect 26236 5842 26292 5854
rect 26348 3554 26404 9436
rect 26460 8260 26516 8270
rect 26460 7588 26516 8204
rect 26460 5906 26516 7532
rect 26796 8146 26852 8158
rect 26796 8094 26798 8146
rect 26850 8094 26852 8146
rect 26796 7476 26852 8094
rect 26796 7410 26852 7420
rect 26684 7364 26740 7374
rect 26684 7270 26740 7308
rect 26572 7250 26628 7262
rect 26572 7198 26574 7250
rect 26626 7198 26628 7250
rect 26572 7140 26628 7198
rect 26572 7074 26628 7084
rect 26796 7028 26852 7038
rect 26796 6130 26852 6972
rect 26796 6078 26798 6130
rect 26850 6078 26852 6130
rect 26796 6066 26852 6078
rect 26460 5854 26462 5906
rect 26514 5854 26516 5906
rect 26460 5842 26516 5854
rect 26460 5348 26516 5358
rect 26460 4450 26516 5292
rect 26796 5236 26852 5246
rect 26908 5236 26964 11732
rect 27020 7924 27076 12124
rect 27244 11844 27300 11854
rect 27132 11170 27188 11182
rect 27132 11118 27134 11170
rect 27186 11118 27188 11170
rect 27132 8484 27188 11118
rect 27132 8418 27188 8428
rect 27020 7858 27076 7868
rect 27132 7474 27188 7486
rect 27132 7422 27134 7474
rect 27186 7422 27188 7474
rect 27132 7252 27188 7422
rect 27132 7186 27188 7196
rect 26796 5234 26964 5236
rect 26796 5182 26798 5234
rect 26850 5182 26964 5234
rect 26796 5180 26964 5182
rect 26796 5170 26852 5180
rect 26460 4398 26462 4450
rect 26514 4398 26516 4450
rect 26460 4386 26516 4398
rect 26684 5012 26740 5022
rect 26348 3502 26350 3554
rect 26402 3502 26404 3554
rect 26348 3490 26404 3502
rect 25452 3378 25508 3388
rect 25788 3332 26068 3388
rect 25788 2772 25844 3332
rect 25788 2706 25844 2716
rect 26684 800 26740 4956
rect 27244 3554 27300 11788
rect 27356 11396 27412 12798
rect 27468 12852 27524 12862
rect 27468 12758 27524 12796
rect 27468 12292 27524 12302
rect 27468 12198 27524 12236
rect 27580 11508 27636 13692
rect 27692 12852 27748 15148
rect 27692 12786 27748 12796
rect 27804 11956 27860 15820
rect 28252 15874 28308 15886
rect 28252 15822 28254 15874
rect 28306 15822 28308 15874
rect 28252 15428 28308 15822
rect 28252 15362 28308 15372
rect 28812 15874 28868 15886
rect 28812 15822 28814 15874
rect 28866 15822 28868 15874
rect 28028 15316 28084 15326
rect 28084 15260 28196 15316
rect 28028 15222 28084 15260
rect 28140 15148 28196 15260
rect 28588 15202 28644 15214
rect 28588 15150 28590 15202
rect 28642 15150 28644 15202
rect 28140 15092 28420 15148
rect 28028 14644 28084 14654
rect 28028 14550 28084 14588
rect 28140 13972 28196 13982
rect 28140 13878 28196 13916
rect 27916 13746 27972 13758
rect 28252 13748 28308 13758
rect 27916 13694 27918 13746
rect 27970 13694 27972 13746
rect 27916 12964 27972 13694
rect 28140 13746 28308 13748
rect 28140 13694 28254 13746
rect 28306 13694 28308 13746
rect 28140 13692 28308 13694
rect 28140 13300 28196 13692
rect 28252 13682 28308 13692
rect 28364 13524 28420 15092
rect 28140 13234 28196 13244
rect 28252 13468 28420 13524
rect 28476 14306 28532 14318
rect 28476 14254 28478 14306
rect 28530 14254 28532 14306
rect 27916 12898 27972 12908
rect 28252 12850 28308 13468
rect 28476 13300 28532 14254
rect 28476 13234 28532 13244
rect 28588 13524 28644 15150
rect 28812 14308 28868 15822
rect 30716 15540 30772 15550
rect 30716 15446 30772 15484
rect 30044 15428 30100 15438
rect 29820 15316 29876 15326
rect 29820 15222 29876 15260
rect 28812 14242 28868 14252
rect 28924 15204 28980 15214
rect 28812 13748 28868 13758
rect 28812 13634 28868 13692
rect 28812 13582 28814 13634
rect 28866 13582 28868 13634
rect 28812 13524 28868 13582
rect 28588 13468 28868 13524
rect 28924 13522 28980 15148
rect 29036 15202 29092 15214
rect 29036 15150 29038 15202
rect 29090 15150 29092 15202
rect 29036 13972 29092 15150
rect 29484 15202 29540 15214
rect 29484 15150 29486 15202
rect 29538 15150 29540 15202
rect 29484 15148 29540 15150
rect 29036 13906 29092 13916
rect 29372 15092 29540 15148
rect 29372 13636 29428 15092
rect 29372 13542 29428 13580
rect 29484 14308 29540 14318
rect 28924 13470 28926 13522
rect 28978 13470 28980 13522
rect 28588 13076 28644 13468
rect 28252 12798 28254 12850
rect 28306 12798 28308 12850
rect 28252 12786 28308 12798
rect 28364 13020 28644 13076
rect 28364 12850 28420 13020
rect 28364 12798 28366 12850
rect 28418 12798 28420 12850
rect 27804 11890 27860 11900
rect 28028 12738 28084 12750
rect 28028 12686 28030 12738
rect 28082 12686 28084 12738
rect 27916 11508 27972 11518
rect 27580 11506 27972 11508
rect 27580 11454 27918 11506
rect 27970 11454 27972 11506
rect 27580 11452 27972 11454
rect 27916 11442 27972 11452
rect 27356 11330 27412 11340
rect 27468 11282 27524 11294
rect 27468 11230 27470 11282
rect 27522 11230 27524 11282
rect 27356 11172 27412 11182
rect 27356 11078 27412 11116
rect 27468 11060 27524 11230
rect 27468 10724 27524 11004
rect 27468 10658 27524 10668
rect 27356 10500 27412 10510
rect 27356 10050 27412 10444
rect 27356 9998 27358 10050
rect 27410 9998 27412 10050
rect 27356 9986 27412 9998
rect 27580 10052 27636 10062
rect 27804 10052 27860 10062
rect 27636 9996 27748 10052
rect 27580 9986 27636 9996
rect 27468 9940 27524 9950
rect 27468 9846 27524 9884
rect 27692 9938 27748 9996
rect 27804 9958 27860 9996
rect 27692 9886 27694 9938
rect 27746 9886 27748 9938
rect 27692 9380 27748 9886
rect 27692 9314 27748 9324
rect 27692 9156 27748 9166
rect 27580 7700 27636 7710
rect 27468 7644 27580 7700
rect 27468 5906 27524 7644
rect 27580 7606 27636 7644
rect 27692 7698 27748 9100
rect 27804 8932 27860 8942
rect 27804 8838 27860 8876
rect 27692 7646 27694 7698
rect 27746 7646 27748 7698
rect 27692 7634 27748 7646
rect 27804 8260 27860 8270
rect 27804 7698 27860 8204
rect 27804 7646 27806 7698
rect 27858 7646 27860 7698
rect 27804 7634 27860 7646
rect 27468 5854 27470 5906
rect 27522 5854 27524 5906
rect 27468 5842 27524 5854
rect 27692 6468 27748 6478
rect 27692 5906 27748 6412
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 27692 5842 27748 5854
rect 28028 5906 28084 12686
rect 28364 12516 28420 12798
rect 28364 12450 28420 12460
rect 28812 12738 28868 12750
rect 28812 12686 28814 12738
rect 28866 12686 28868 12738
rect 28812 12516 28868 12686
rect 28812 12450 28868 12460
rect 28812 12292 28868 12302
rect 28364 12068 28420 12078
rect 28252 11956 28308 11966
rect 28252 8260 28308 11900
rect 28364 11394 28420 12012
rect 28700 11620 28756 11630
rect 28364 11342 28366 11394
rect 28418 11342 28420 11394
rect 28364 11330 28420 11342
rect 28588 11508 28644 11518
rect 28588 11170 28644 11452
rect 28700 11394 28756 11564
rect 28700 11342 28702 11394
rect 28754 11342 28756 11394
rect 28700 11330 28756 11342
rect 28812 11172 28868 12236
rect 28588 11118 28590 11170
rect 28642 11118 28644 11170
rect 28588 10836 28644 11118
rect 28588 10770 28644 10780
rect 28700 11116 28868 11172
rect 28700 10500 28756 11116
rect 28924 10948 28980 13470
rect 29372 11956 29428 11966
rect 28924 10892 29204 10948
rect 28924 10500 28980 10510
rect 28700 10498 28980 10500
rect 28700 10446 28926 10498
rect 28978 10446 28980 10498
rect 28700 10444 28980 10446
rect 28476 9940 28532 9950
rect 28476 9846 28532 9884
rect 28700 9716 28756 10444
rect 28924 10434 28980 10444
rect 29148 10276 29204 10892
rect 28924 10220 29204 10276
rect 29260 10724 29316 10734
rect 28812 9716 28868 9726
rect 28700 9714 28868 9716
rect 28700 9662 28814 9714
rect 28866 9662 28868 9714
rect 28700 9660 28868 9662
rect 28588 9604 28644 9614
rect 28588 9602 28756 9604
rect 28588 9550 28590 9602
rect 28642 9550 28756 9602
rect 28588 9548 28756 9550
rect 28588 9538 28644 9548
rect 28588 9044 28644 9054
rect 28588 8950 28644 8988
rect 28700 8820 28756 9548
rect 28252 8194 28308 8204
rect 28588 8764 28756 8820
rect 28588 8372 28644 8764
rect 28588 8036 28644 8316
rect 28364 7980 28644 8036
rect 28700 8034 28756 8046
rect 28700 7982 28702 8034
rect 28754 7982 28756 8034
rect 28252 6804 28308 6814
rect 28252 6690 28308 6748
rect 28252 6638 28254 6690
rect 28306 6638 28308 6690
rect 28252 6626 28308 6638
rect 28364 6132 28420 7980
rect 28476 7476 28532 7486
rect 28532 7420 28644 7476
rect 28476 7344 28532 7420
rect 28588 6468 28644 7420
rect 28700 6914 28756 7982
rect 28700 6862 28702 6914
rect 28754 6862 28756 6914
rect 28700 6850 28756 6862
rect 28700 6468 28756 6478
rect 28588 6466 28756 6468
rect 28588 6414 28702 6466
rect 28754 6414 28756 6466
rect 28588 6412 28756 6414
rect 28476 6132 28532 6142
rect 28364 6130 28532 6132
rect 28364 6078 28478 6130
rect 28530 6078 28532 6130
rect 28364 6076 28532 6078
rect 28476 6066 28532 6076
rect 28588 6020 28644 6030
rect 28588 5926 28644 5964
rect 28028 5854 28030 5906
rect 28082 5854 28084 5906
rect 28028 5842 28084 5854
rect 27804 5794 27860 5806
rect 27804 5742 27806 5794
rect 27858 5742 27860 5794
rect 27804 5236 27860 5742
rect 27804 5170 27860 5180
rect 28476 5122 28532 5134
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 27468 5012 27524 5022
rect 27468 4918 27524 4956
rect 28476 4564 28532 5070
rect 28700 5124 28756 6412
rect 28700 5058 28756 5068
rect 28476 4498 28532 4508
rect 28812 4340 28868 9660
rect 28924 7140 28980 10220
rect 29260 9268 29316 10668
rect 28924 7074 28980 7084
rect 29036 9212 29316 9268
rect 28924 6914 28980 6926
rect 28924 6862 28926 6914
rect 28978 6862 28980 6914
rect 28924 6244 28980 6862
rect 28924 6178 28980 6188
rect 29036 6020 29092 9212
rect 29260 9042 29316 9054
rect 29260 8990 29262 9042
rect 29314 8990 29316 9042
rect 29148 8820 29204 8830
rect 29148 7586 29204 8764
rect 29148 7534 29150 7586
rect 29202 7534 29204 7586
rect 29148 7522 29204 7534
rect 29260 7028 29316 8990
rect 29260 6962 29316 6972
rect 29372 6804 29428 11900
rect 29484 11284 29540 14252
rect 29596 14306 29652 14318
rect 29596 14254 29598 14306
rect 29650 14254 29652 14306
rect 29596 13522 29652 14254
rect 29932 14308 29988 14318
rect 29932 14214 29988 14252
rect 29820 13748 29876 13758
rect 29820 13654 29876 13692
rect 29596 13470 29598 13522
rect 29650 13470 29652 13522
rect 29596 12850 29652 13470
rect 29596 12798 29598 12850
rect 29650 12798 29652 12850
rect 29596 12516 29652 12798
rect 29708 12740 29764 12750
rect 29708 12738 29876 12740
rect 29708 12686 29710 12738
rect 29762 12686 29876 12738
rect 29708 12684 29876 12686
rect 29708 12674 29764 12684
rect 29596 12460 29764 12516
rect 29596 12066 29652 12078
rect 29596 12014 29598 12066
rect 29650 12014 29652 12066
rect 29596 11620 29652 12014
rect 29596 11554 29652 11564
rect 29596 11284 29652 11294
rect 29484 11282 29652 11284
rect 29484 11230 29598 11282
rect 29650 11230 29652 11282
rect 29484 11228 29652 11230
rect 29484 11060 29540 11228
rect 29596 11218 29652 11228
rect 29484 10164 29540 11004
rect 29708 11170 29764 12460
rect 29708 11118 29710 11170
rect 29762 11118 29764 11170
rect 29484 10098 29540 10108
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29036 5954 29092 5964
rect 29260 6748 29428 6804
rect 29484 9154 29540 9166
rect 29484 9102 29486 9154
rect 29538 9102 29540 9154
rect 29260 5906 29316 6748
rect 29372 6132 29428 6142
rect 29372 6038 29428 6076
rect 29260 5854 29262 5906
rect 29314 5854 29316 5906
rect 29260 5842 29316 5854
rect 29036 5124 29092 5134
rect 29036 4562 29092 5068
rect 29036 4510 29038 4562
rect 29090 4510 29092 4562
rect 29036 4498 29092 4510
rect 28812 4274 28868 4284
rect 28588 4228 28644 4238
rect 28588 4134 28644 4172
rect 27804 3668 27860 3678
rect 27804 3574 27860 3612
rect 28028 3668 28084 3678
rect 27244 3502 27246 3554
rect 27298 3502 27300 3554
rect 27244 3490 27300 3502
rect 28028 800 28084 3612
rect 29484 3554 29540 9102
rect 29596 9044 29652 10558
rect 29708 10388 29764 11118
rect 29820 11620 29876 12684
rect 29820 11172 29876 11564
rect 29932 11396 29988 11406
rect 30044 11396 30100 15372
rect 31164 15428 31220 15438
rect 31164 15334 31220 15372
rect 31948 15316 32004 15326
rect 30380 15204 30436 15214
rect 30380 15110 30436 15148
rect 31724 15202 31780 15214
rect 31724 15150 31726 15202
rect 31778 15150 31780 15202
rect 30380 14308 30436 14318
rect 30940 14308 30996 14318
rect 30380 14306 30548 14308
rect 30380 14254 30382 14306
rect 30434 14254 30548 14306
rect 30380 14252 30548 14254
rect 30380 14242 30436 14252
rect 30268 13634 30324 13646
rect 30268 13582 30270 13634
rect 30322 13582 30324 13634
rect 30268 13522 30324 13582
rect 30268 13470 30270 13522
rect 30322 13470 30324 13522
rect 30268 13458 30324 13470
rect 30268 12852 30324 12890
rect 30268 12786 30324 12796
rect 30380 12738 30436 12750
rect 30380 12686 30382 12738
rect 30434 12686 30436 12738
rect 30268 12628 30324 12638
rect 30268 12290 30324 12572
rect 30268 12238 30270 12290
rect 30322 12238 30324 12290
rect 30268 12226 30324 12238
rect 30156 12180 30212 12190
rect 30156 12086 30212 12124
rect 30380 11844 30436 12686
rect 30492 12068 30548 14252
rect 30940 14214 30996 14252
rect 31612 14308 31668 14318
rect 30716 13634 30772 13646
rect 30716 13582 30718 13634
rect 30770 13582 30772 13634
rect 30716 12740 30772 13582
rect 31164 13636 31220 13646
rect 31164 13542 31220 13580
rect 30716 12674 30772 12684
rect 30940 12850 30996 12862
rect 30940 12798 30942 12850
rect 30994 12798 30996 12850
rect 30940 12292 30996 12798
rect 31276 12852 31332 12862
rect 30716 12236 30996 12292
rect 31052 12738 31108 12750
rect 31052 12686 31054 12738
rect 31106 12686 31108 12738
rect 30604 12068 30660 12078
rect 30492 12012 30604 12068
rect 30380 11778 30436 11788
rect 29988 11340 30100 11396
rect 30604 11394 30660 12012
rect 30604 11342 30606 11394
rect 30658 11342 30660 11394
rect 29932 11264 29988 11340
rect 30604 11330 30660 11342
rect 29876 11116 29988 11172
rect 29820 11040 29876 11116
rect 29708 10322 29764 10332
rect 29596 8978 29652 8988
rect 29708 10164 29764 10174
rect 29596 7028 29652 7038
rect 29596 6914 29652 6972
rect 29596 6862 29598 6914
rect 29650 6862 29652 6914
rect 29596 6850 29652 6862
rect 29596 6244 29652 6254
rect 29708 6244 29764 10108
rect 29820 9826 29876 9838
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 29820 9268 29876 9774
rect 29820 9202 29876 9212
rect 29932 9156 29988 11116
rect 30268 11170 30324 11182
rect 30268 11118 30270 11170
rect 30322 11118 30324 11170
rect 30268 10724 30324 11118
rect 30268 10658 30324 10668
rect 30380 11172 30436 11182
rect 30268 10498 30324 10510
rect 30268 10446 30270 10498
rect 30322 10446 30324 10498
rect 30156 9940 30212 9950
rect 30268 9940 30324 10446
rect 30156 9938 30324 9940
rect 30156 9886 30158 9938
rect 30210 9886 30324 9938
rect 30156 9884 30324 9886
rect 30156 9874 30212 9884
rect 30044 9828 30100 9838
rect 30044 9734 30100 9772
rect 30380 9826 30436 11116
rect 30380 9774 30382 9826
rect 30434 9774 30436 9826
rect 30380 9762 30436 9774
rect 30492 11170 30548 11182
rect 30492 11118 30494 11170
rect 30546 11118 30548 11170
rect 30380 9492 30436 9502
rect 30268 9156 30324 9166
rect 29932 9100 30212 9156
rect 30044 8818 30100 8830
rect 30044 8766 30046 8818
rect 30098 8766 30100 8818
rect 30044 8372 30100 8766
rect 30044 8306 30100 8316
rect 29820 8258 29876 8270
rect 29820 8206 29822 8258
rect 29874 8206 29876 8258
rect 29820 7252 29876 8206
rect 29820 7186 29876 7196
rect 29932 8260 29988 8270
rect 29932 7700 29988 8204
rect 30156 7812 30212 9100
rect 30268 9062 30324 9100
rect 30268 8932 30324 8942
rect 30268 8838 30324 8876
rect 30380 8258 30436 9436
rect 30380 8206 30382 8258
rect 30434 8206 30436 8258
rect 30380 8194 30436 8206
rect 30492 8260 30548 11118
rect 30716 11172 30772 12236
rect 30940 12068 30996 12078
rect 30940 11974 30996 12012
rect 30828 11956 30884 11966
rect 30828 11862 30884 11900
rect 31052 11508 31108 12686
rect 31052 11442 31108 11452
rect 31052 11284 31108 11294
rect 31052 11190 31108 11228
rect 30716 11106 30772 11116
rect 30492 8194 30548 8204
rect 30604 10052 30660 10062
rect 30268 8036 30324 8046
rect 30268 7942 30324 7980
rect 30492 8034 30548 8046
rect 30492 7982 30494 8034
rect 30546 7982 30548 8034
rect 30156 7756 30436 7812
rect 29932 6914 29988 7644
rect 29932 6862 29934 6914
rect 29986 6862 29988 6914
rect 29932 6850 29988 6862
rect 29820 6468 29876 6478
rect 29820 6374 29876 6412
rect 30380 6356 30436 7756
rect 30492 7364 30548 7982
rect 30604 8036 30660 9996
rect 31052 9828 31108 9838
rect 30940 9492 30996 9502
rect 30940 9042 30996 9436
rect 30940 8990 30942 9042
rect 30994 8990 30996 9042
rect 30940 8978 30996 8990
rect 31052 8932 31108 9772
rect 31164 9716 31220 9726
rect 31164 9622 31220 9660
rect 31276 9492 31332 12796
rect 31612 12740 31668 14252
rect 31724 13860 31780 15150
rect 31948 14754 32004 15260
rect 32172 15204 32228 15214
rect 32620 15204 32676 15214
rect 32172 15202 32340 15204
rect 32172 15150 32174 15202
rect 32226 15150 32340 15202
rect 32172 15148 32340 15150
rect 32172 15138 32228 15148
rect 31948 14702 31950 14754
rect 32002 14702 32004 14754
rect 31948 14690 32004 14702
rect 32060 14306 32116 14318
rect 32060 14254 32062 14306
rect 32114 14254 32116 14306
rect 31724 13794 31780 13804
rect 31948 13972 32004 13982
rect 31724 13636 31780 13646
rect 31724 13634 31892 13636
rect 31724 13582 31726 13634
rect 31778 13582 31892 13634
rect 31724 13580 31892 13582
rect 31724 13570 31780 13580
rect 31388 12738 31668 12740
rect 31388 12686 31614 12738
rect 31666 12686 31668 12738
rect 31388 12684 31668 12686
rect 31388 9828 31444 12684
rect 31612 12674 31668 12684
rect 31724 12850 31780 12862
rect 31724 12798 31726 12850
rect 31778 12798 31780 12850
rect 31612 12066 31668 12078
rect 31612 12014 31614 12066
rect 31666 12014 31668 12066
rect 31500 11956 31556 11966
rect 31500 11862 31556 11900
rect 31388 9762 31444 9772
rect 31500 11508 31556 11518
rect 30940 8820 30996 8830
rect 30940 8726 30996 8764
rect 31052 8596 31108 8876
rect 30604 7970 30660 7980
rect 30716 8540 31108 8596
rect 31164 9436 31332 9492
rect 31500 9714 31556 11452
rect 31500 9662 31502 9714
rect 31554 9662 31556 9714
rect 30492 7298 30548 7308
rect 30604 6692 30660 6702
rect 30604 6598 30660 6636
rect 30492 6580 30548 6590
rect 30492 6486 30548 6524
rect 30380 6300 30548 6356
rect 29652 6188 29764 6244
rect 29596 6130 29652 6188
rect 29596 6078 29598 6130
rect 29650 6078 29652 6130
rect 29596 6066 29652 6078
rect 29932 6020 29988 6030
rect 29932 5926 29988 5964
rect 29820 5908 29876 5918
rect 29820 5814 29876 5852
rect 30380 5908 30436 5918
rect 30380 5814 30436 5852
rect 30492 5906 30548 6300
rect 30492 5854 30494 5906
rect 30546 5854 30548 5906
rect 30492 5842 30548 5854
rect 30716 5906 30772 8540
rect 31052 8372 31108 8382
rect 30828 8370 31108 8372
rect 30828 8318 31054 8370
rect 31106 8318 31108 8370
rect 30828 8316 31108 8318
rect 30828 7028 30884 8316
rect 31052 8306 31108 8316
rect 31164 8370 31220 9436
rect 31500 9380 31556 9662
rect 31276 9324 31556 9380
rect 31612 11396 31668 12014
rect 31724 11732 31780 12798
rect 31836 12068 31892 13580
rect 31836 12002 31892 12012
rect 31948 11844 32004 13916
rect 31724 11666 31780 11676
rect 31836 11788 32004 11844
rect 32060 12066 32116 14254
rect 32284 14084 32340 15148
rect 32620 15110 32676 15148
rect 33740 15204 33796 15214
rect 33516 14754 33572 14766
rect 33516 14702 33518 14754
rect 33570 14702 33572 14754
rect 32844 14532 32900 14542
rect 32396 14308 32452 14318
rect 32396 14214 32452 14252
rect 32844 14306 32900 14476
rect 33292 14420 33348 14430
rect 33292 14326 33348 14364
rect 32844 14254 32846 14306
rect 32898 14254 32900 14306
rect 32284 14028 32452 14084
rect 32172 13972 32228 13982
rect 32172 13878 32228 13916
rect 32284 13860 32340 13870
rect 32172 13188 32228 13198
rect 32172 12292 32228 13132
rect 32172 12226 32228 12236
rect 32284 12964 32340 13804
rect 32396 13188 32452 14028
rect 32620 13636 32676 13646
rect 32620 13542 32676 13580
rect 32844 13188 32900 14254
rect 33404 13636 33460 13646
rect 32844 13132 33236 13188
rect 32396 13122 32452 13132
rect 32844 12964 32900 12974
rect 32284 12962 32900 12964
rect 32284 12910 32846 12962
rect 32898 12910 32900 12962
rect 32284 12908 32900 12910
rect 32284 12850 32340 12908
rect 32844 12898 32900 12908
rect 32284 12798 32286 12850
rect 32338 12798 32340 12850
rect 32060 12014 32062 12066
rect 32114 12014 32116 12066
rect 31724 11396 31780 11406
rect 31612 11394 31780 11396
rect 31612 11342 31726 11394
rect 31778 11342 31780 11394
rect 31612 11340 31780 11342
rect 31276 9154 31332 9324
rect 31276 9102 31278 9154
rect 31330 9102 31332 9154
rect 31276 9090 31332 9102
rect 31164 8318 31166 8370
rect 31218 8318 31220 8370
rect 30828 6962 30884 6972
rect 30940 8148 30996 8158
rect 30716 5854 30718 5906
rect 30770 5854 30772 5906
rect 30716 5842 30772 5854
rect 30940 5906 30996 8092
rect 31164 7140 31220 8318
rect 31388 8260 31444 8270
rect 31388 8166 31444 8204
rect 31276 7364 31332 7374
rect 31612 7364 31668 11340
rect 31724 11330 31780 11340
rect 31836 11282 31892 11788
rect 32060 11620 32116 12014
rect 32060 11554 32116 11564
rect 31836 11230 31838 11282
rect 31890 11230 31892 11282
rect 31836 10724 31892 11230
rect 32060 11172 32116 11182
rect 32060 11078 32116 11116
rect 31724 10668 31892 10724
rect 31724 10052 31780 10668
rect 31724 9986 31780 9996
rect 31836 10500 31892 10510
rect 31836 9826 31892 10444
rect 31836 9774 31838 9826
rect 31890 9774 31892 9826
rect 31836 9762 31892 9774
rect 31836 9604 31892 9614
rect 31836 9602 32004 9604
rect 31836 9550 31838 9602
rect 31890 9550 32004 9602
rect 31836 9548 32004 9550
rect 31836 9538 31892 9548
rect 31724 9044 31780 9054
rect 31724 8372 31780 8988
rect 31836 8932 31892 8942
rect 31836 8838 31892 8876
rect 31836 8372 31892 8382
rect 31724 8370 31892 8372
rect 31724 8318 31838 8370
rect 31890 8318 31892 8370
rect 31724 8316 31892 8318
rect 31836 8306 31892 8316
rect 31948 7924 32004 9548
rect 32060 9492 32116 9502
rect 32060 9266 32116 9436
rect 32060 9214 32062 9266
rect 32114 9214 32116 9266
rect 32060 9202 32116 9214
rect 32284 9044 32340 12798
rect 32396 12740 32452 12750
rect 32396 12738 33124 12740
rect 32396 12686 32398 12738
rect 32450 12686 33124 12738
rect 32396 12684 33124 12686
rect 32396 12674 32452 12684
rect 32956 12516 33012 12526
rect 32732 12292 32788 12302
rect 32732 12198 32788 12236
rect 32844 12180 32900 12190
rect 32844 12086 32900 12124
rect 32732 11954 32788 11966
rect 32732 11902 32734 11954
rect 32786 11902 32788 11954
rect 32396 11732 32452 11742
rect 32396 11284 32452 11676
rect 32620 11508 32676 11518
rect 32508 11284 32564 11294
rect 32396 11282 32564 11284
rect 32396 11230 32510 11282
rect 32562 11230 32564 11282
rect 32396 11228 32564 11230
rect 32396 10500 32452 11228
rect 32508 11218 32564 11228
rect 32620 11282 32676 11452
rect 32620 11230 32622 11282
rect 32674 11230 32676 11282
rect 32620 11218 32676 11230
rect 32396 10406 32452 10444
rect 32060 8988 32340 9044
rect 32508 9826 32564 9838
rect 32508 9774 32510 9826
rect 32562 9774 32564 9826
rect 32508 9044 32564 9774
rect 32620 9380 32676 9390
rect 32620 9266 32676 9324
rect 32620 9214 32622 9266
rect 32674 9214 32676 9266
rect 32620 9202 32676 9214
rect 32060 8596 32116 8988
rect 32508 8978 32564 8988
rect 32172 8820 32228 8830
rect 32396 8820 32452 8830
rect 32172 8818 32452 8820
rect 32172 8766 32174 8818
rect 32226 8766 32398 8818
rect 32450 8766 32452 8818
rect 32172 8764 32452 8766
rect 32172 8754 32228 8764
rect 32396 8754 32452 8764
rect 32060 8540 32228 8596
rect 31948 7586 32004 7868
rect 31948 7534 31950 7586
rect 32002 7534 32004 7586
rect 31948 7522 32004 7534
rect 31332 7308 31668 7364
rect 32060 7362 32116 7374
rect 32060 7310 32062 7362
rect 32114 7310 32116 7362
rect 31276 7232 31332 7308
rect 31052 7084 31220 7140
rect 31052 6132 31108 7084
rect 31052 6066 31108 6076
rect 31164 6916 31220 6926
rect 31164 6690 31220 6860
rect 31948 6804 32004 6814
rect 32060 6804 32116 7310
rect 31948 6802 32116 6804
rect 31948 6750 31950 6802
rect 32002 6750 32116 6802
rect 31948 6748 32116 6750
rect 31948 6738 32004 6748
rect 31164 6638 31166 6690
rect 31218 6638 31220 6690
rect 30940 5854 30942 5906
rect 30994 5854 30996 5906
rect 30940 5842 30996 5854
rect 30716 5236 30772 5246
rect 30716 5142 30772 5180
rect 29932 5124 29988 5134
rect 29932 5030 29988 5068
rect 31164 5124 31220 6638
rect 32172 6132 32228 8540
rect 32508 8372 32564 8382
rect 32508 8260 32564 8316
rect 32284 8258 32564 8260
rect 32284 8206 32510 8258
rect 32562 8206 32564 8258
rect 32284 8204 32564 8206
rect 32284 7586 32340 8204
rect 32508 8194 32564 8204
rect 32732 8260 32788 11902
rect 32844 11172 32900 11182
rect 32844 11078 32900 11116
rect 32844 10836 32900 10846
rect 32956 10836 33012 12460
rect 32844 10834 33012 10836
rect 32844 10782 32846 10834
rect 32898 10782 33012 10834
rect 32844 10780 33012 10782
rect 32844 10770 32900 10780
rect 33068 9604 33124 12684
rect 33180 11956 33236 13132
rect 33292 12738 33348 12750
rect 33292 12686 33294 12738
rect 33346 12686 33348 12738
rect 33292 12180 33348 12686
rect 33404 12404 33460 13580
rect 33516 13634 33572 14702
rect 33516 13582 33518 13634
rect 33570 13582 33572 13634
rect 33516 13186 33572 13582
rect 33516 13134 33518 13186
rect 33570 13134 33572 13186
rect 33516 13122 33572 13134
rect 33628 13522 33684 13534
rect 33628 13470 33630 13522
rect 33682 13470 33684 13522
rect 33516 12404 33572 12414
rect 33404 12402 33572 12404
rect 33404 12350 33518 12402
rect 33570 12350 33572 12402
rect 33404 12348 33572 12350
rect 33292 12114 33348 12124
rect 33180 11900 33348 11956
rect 33180 11396 33236 11406
rect 33180 11302 33236 11340
rect 33292 10948 33348 11900
rect 33516 11954 33572 12348
rect 33516 11902 33518 11954
rect 33570 11902 33572 11954
rect 33516 11890 33572 11902
rect 33628 11396 33684 13470
rect 33740 13074 33796 15148
rect 33740 13022 33742 13074
rect 33794 13022 33796 13074
rect 33740 13010 33796 13022
rect 33852 14306 33908 14318
rect 33852 14254 33854 14306
rect 33906 14254 33908 14306
rect 33852 12180 33908 14254
rect 34300 14306 34356 16156
rect 36540 15428 36596 15438
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34300 14254 34302 14306
rect 34354 14254 34356 14306
rect 34076 13634 34132 13646
rect 34076 13582 34078 13634
rect 34130 13582 34132 13634
rect 33964 12292 34020 12302
rect 33964 12198 34020 12236
rect 33516 11172 33572 11182
rect 33068 9538 33124 9548
rect 33180 10892 33348 10948
rect 33404 10948 33460 10958
rect 32732 8194 32788 8204
rect 32956 9044 33012 9054
rect 32284 7534 32286 7586
rect 32338 7534 32340 7586
rect 32284 7522 32340 7534
rect 32396 8036 32452 8046
rect 32172 6066 32228 6076
rect 31500 6020 31556 6030
rect 31500 5926 31556 5964
rect 31836 6020 31892 6030
rect 31836 5926 31892 5964
rect 32060 5906 32116 5918
rect 32060 5854 32062 5906
rect 32114 5854 32116 5906
rect 31612 5794 31668 5806
rect 31612 5742 31614 5794
rect 31666 5742 31668 5794
rect 31164 5058 31220 5068
rect 31388 5348 31444 5358
rect 30828 4452 30884 4462
rect 30828 4338 30884 4396
rect 30828 4286 30830 4338
rect 30882 4286 30884 4338
rect 30828 4274 30884 4286
rect 31388 4338 31444 5292
rect 31612 5236 31668 5742
rect 32060 5796 32116 5854
rect 32060 5730 32116 5740
rect 32284 5908 32340 5918
rect 31612 5170 31668 5180
rect 31388 4286 31390 4338
rect 31442 4286 31444 4338
rect 31388 4274 31444 4286
rect 31612 4340 31668 4350
rect 31612 4246 31668 4284
rect 31948 4340 32004 4350
rect 31948 4246 32004 4284
rect 29484 3502 29486 3554
rect 29538 3502 29540 3554
rect 29484 3490 29540 3502
rect 29708 4226 29764 4238
rect 29708 4174 29710 4226
rect 29762 4174 29764 4226
rect 29708 3388 29764 4174
rect 29932 3668 29988 3678
rect 29932 3574 29988 3612
rect 32172 3668 32228 3678
rect 31164 3442 31220 3454
rect 31164 3390 31166 3442
rect 31218 3390 31220 3442
rect 31164 3388 31220 3390
rect 29596 3332 29764 3388
rect 30716 3332 31220 3388
rect 29596 980 29652 3332
rect 29372 924 29652 980
rect 29372 800 29428 924
rect 30716 800 30772 3332
rect 32172 1764 32228 3612
rect 32284 3554 32340 5852
rect 32396 4340 32452 7980
rect 32620 8034 32676 8046
rect 32620 7982 32622 8034
rect 32674 7982 32676 8034
rect 32508 7588 32564 7598
rect 32620 7588 32676 7982
rect 32732 8034 32788 8046
rect 32732 7982 32734 8034
rect 32786 7982 32788 8034
rect 32732 7924 32788 7982
rect 32732 7858 32788 7868
rect 32956 8034 33012 8988
rect 32956 7982 32958 8034
rect 33010 7982 33012 8034
rect 32508 7586 32676 7588
rect 32508 7534 32510 7586
rect 32562 7534 32676 7586
rect 32508 7532 32676 7534
rect 32508 7522 32564 7532
rect 32956 7252 33012 7982
rect 32956 7186 33012 7196
rect 33068 8818 33124 8830
rect 33068 8766 33070 8818
rect 33122 8766 33124 8818
rect 32956 7028 33012 7038
rect 32732 6356 32788 6366
rect 32732 6018 32788 6300
rect 32732 5966 32734 6018
rect 32786 5966 32788 6018
rect 32508 5906 32564 5918
rect 32508 5854 32510 5906
rect 32562 5854 32564 5906
rect 32508 5124 32564 5854
rect 32732 5684 32788 5966
rect 32844 6244 32900 6254
rect 32844 6018 32900 6188
rect 32844 5966 32846 6018
rect 32898 5966 32900 6018
rect 32844 5954 32900 5966
rect 32732 5618 32788 5628
rect 32844 5236 32900 5246
rect 32844 5142 32900 5180
rect 32508 5058 32564 5068
rect 32732 4564 32788 4574
rect 32732 4470 32788 4508
rect 32844 4452 32900 4462
rect 32956 4452 33012 6972
rect 32844 4450 33012 4452
rect 32844 4398 32846 4450
rect 32898 4398 33012 4450
rect 32844 4396 33012 4398
rect 32844 4386 32900 4396
rect 32508 4340 32564 4350
rect 32396 4338 32564 4340
rect 32396 4286 32510 4338
rect 32562 4286 32564 4338
rect 32396 4284 32564 4286
rect 32508 4274 32564 4284
rect 32284 3502 32286 3554
rect 32338 3502 32340 3554
rect 32284 3490 32340 3502
rect 33068 3556 33124 8766
rect 33180 6356 33236 10892
rect 33292 9940 33348 9950
rect 33292 9846 33348 9884
rect 33180 6290 33236 6300
rect 33404 5348 33460 10892
rect 33516 10612 33572 11116
rect 33628 10948 33684 11340
rect 33628 10882 33684 10892
rect 33740 12124 33908 12180
rect 34076 12180 34132 13582
rect 34188 12738 34244 12750
rect 34188 12686 34190 12738
rect 34242 12686 34244 12738
rect 34188 12516 34244 12686
rect 34300 12740 34356 14254
rect 34748 13972 34804 13982
rect 34300 12674 34356 12684
rect 34524 13634 34580 13646
rect 34524 13582 34526 13634
rect 34578 13582 34580 13634
rect 34188 12450 34244 12460
rect 34076 12124 34356 12180
rect 33740 10724 33796 12124
rect 33852 11954 33908 11966
rect 33852 11902 33854 11954
rect 33906 11902 33908 11954
rect 33852 11394 33908 11902
rect 33852 11342 33854 11394
rect 33906 11342 33908 11394
rect 33852 11330 33908 11342
rect 33964 11956 34020 11966
rect 33740 10668 33908 10724
rect 33516 10610 33684 10612
rect 33516 10558 33518 10610
rect 33570 10558 33684 10610
rect 33516 10556 33684 10558
rect 33516 10546 33572 10556
rect 33516 9268 33572 9278
rect 33628 9268 33684 10556
rect 33740 10498 33796 10510
rect 33740 10446 33742 10498
rect 33794 10446 33796 10498
rect 33740 9940 33796 10446
rect 33740 9874 33796 9884
rect 33852 9828 33908 10668
rect 33852 9762 33908 9772
rect 33964 10722 34020 11900
rect 33964 10670 33966 10722
rect 34018 10670 34020 10722
rect 33740 9268 33796 9278
rect 33628 9266 33796 9268
rect 33628 9214 33742 9266
rect 33794 9214 33796 9266
rect 33628 9212 33796 9214
rect 33516 9174 33572 9212
rect 33740 9202 33796 9212
rect 33852 9044 33908 9054
rect 33852 8950 33908 8988
rect 33628 8708 33684 8718
rect 33628 7586 33684 8652
rect 33964 8708 34020 10670
rect 34188 10612 34244 10622
rect 34188 10518 34244 10556
rect 33964 8642 34020 8652
rect 34188 9828 34244 9838
rect 33740 8260 33796 8270
rect 33740 8036 33796 8204
rect 33964 8148 34020 8158
rect 33964 8054 34020 8092
rect 33740 7942 33796 7980
rect 33852 8034 33908 8046
rect 33852 7982 33854 8034
rect 33906 7982 33908 8034
rect 33852 7812 33908 7982
rect 34076 8036 34132 8046
rect 33628 7534 33630 7586
rect 33682 7534 33684 7586
rect 33628 7522 33684 7534
rect 33740 7756 33908 7812
rect 33964 7812 34020 7822
rect 33404 5234 33460 5292
rect 33404 5182 33406 5234
rect 33458 5182 33460 5234
rect 33404 5170 33460 5182
rect 33628 7028 33684 7038
rect 33628 6018 33684 6972
rect 33628 5966 33630 6018
rect 33682 5966 33684 6018
rect 33628 5346 33684 5966
rect 33740 5908 33796 7756
rect 33852 7588 33908 7598
rect 33852 7494 33908 7532
rect 33964 7362 34020 7756
rect 33964 7310 33966 7362
rect 34018 7310 34020 7362
rect 33964 7298 34020 7310
rect 34076 6802 34132 7980
rect 34188 7028 34244 9772
rect 34300 8372 34356 12124
rect 34412 12066 34468 12078
rect 34412 12014 34414 12066
rect 34466 12014 34468 12066
rect 34412 11954 34468 12014
rect 34412 11902 34414 11954
rect 34466 11902 34468 11954
rect 34412 11890 34468 11902
rect 34524 10836 34580 13582
rect 34748 12964 34804 13916
rect 34860 13634 34916 13646
rect 34860 13582 34862 13634
rect 34914 13582 34916 13634
rect 34860 13522 34916 13582
rect 35420 13636 35476 13646
rect 35420 13634 35812 13636
rect 35420 13582 35422 13634
rect 35474 13582 35812 13634
rect 35420 13580 35812 13582
rect 35420 13570 35476 13580
rect 34860 13470 34862 13522
rect 34914 13470 34916 13522
rect 34860 13458 34916 13470
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34748 12908 34916 12964
rect 34748 12738 34804 12750
rect 34748 12686 34750 12738
rect 34802 12686 34804 12738
rect 34748 12628 34804 12686
rect 34748 12562 34804 12572
rect 34860 12402 34916 12908
rect 35532 12852 35588 12862
rect 35532 12758 35588 12796
rect 35084 12740 35140 12750
rect 35084 12646 35140 12684
rect 34860 12350 34862 12402
rect 34914 12350 34916 12402
rect 34860 12338 34916 12350
rect 34972 12516 35028 12526
rect 34972 11508 35028 12460
rect 35084 12292 35140 12302
rect 35084 11620 35140 12236
rect 35644 12066 35700 12078
rect 35644 12014 35646 12066
rect 35698 12014 35700 12066
rect 35532 11956 35588 11966
rect 35532 11862 35588 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11564 35476 11620
rect 34972 11452 35140 11508
rect 34636 11284 34692 11294
rect 34636 11190 34692 11228
rect 34860 10836 34916 10846
rect 34524 10770 34580 10780
rect 34636 10834 34916 10836
rect 34636 10782 34862 10834
rect 34914 10782 34916 10834
rect 34636 10780 34916 10782
rect 34636 8932 34692 10780
rect 34860 10770 34916 10780
rect 34748 10610 34804 10622
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 34748 9268 34804 10558
rect 34860 10388 34916 10398
rect 34860 10386 35028 10388
rect 34860 10334 34862 10386
rect 34914 10334 35028 10386
rect 34860 10332 35028 10334
rect 34860 10322 34916 10332
rect 34748 9202 34804 9212
rect 34748 9044 34804 9054
rect 34748 9042 34916 9044
rect 34748 8990 34750 9042
rect 34802 8990 34916 9042
rect 34748 8988 34916 8990
rect 34748 8978 34804 8988
rect 34300 7700 34356 8316
rect 34300 7634 34356 7644
rect 34412 8876 34692 8932
rect 34188 6962 34244 6972
rect 34076 6750 34078 6802
rect 34130 6750 34132 6802
rect 34076 6738 34132 6750
rect 34412 6692 34468 8876
rect 34524 8708 34580 8718
rect 34524 8370 34580 8652
rect 34524 8318 34526 8370
rect 34578 8318 34580 8370
rect 34524 8306 34580 8318
rect 34748 8260 34804 8270
rect 34636 8146 34692 8158
rect 34636 8094 34638 8146
rect 34690 8094 34692 8146
rect 34636 7140 34692 8094
rect 34748 8146 34804 8204
rect 34748 8094 34750 8146
rect 34802 8094 34804 8146
rect 34748 8082 34804 8094
rect 34188 6636 34412 6692
rect 33852 6132 33908 6142
rect 33852 6038 33908 6076
rect 34188 6130 34244 6636
rect 34412 6626 34468 6636
rect 34524 7084 34692 7140
rect 34748 7476 34804 7486
rect 34860 7476 34916 8988
rect 34748 7474 34916 7476
rect 34748 7422 34750 7474
rect 34802 7422 34916 7474
rect 34748 7420 34916 7422
rect 34188 6078 34190 6130
rect 34242 6078 34244 6130
rect 34188 6066 34244 6078
rect 33740 5842 33796 5852
rect 34076 6018 34132 6030
rect 34076 5966 34078 6018
rect 34130 5966 34132 6018
rect 33628 5294 33630 5346
rect 33682 5294 33684 5346
rect 33628 5236 33684 5294
rect 34076 5348 34132 5966
rect 34076 5282 34132 5292
rect 33628 5170 33684 5180
rect 33964 5236 34020 5246
rect 33964 5142 34020 5180
rect 33628 4452 33684 4462
rect 33628 4358 33684 4396
rect 33852 4340 33908 4350
rect 33852 4246 33908 4284
rect 34524 4116 34580 7084
rect 34636 6916 34692 6926
rect 34748 6916 34804 7420
rect 34692 6860 34804 6916
rect 34860 7252 34916 7262
rect 34636 5906 34692 6860
rect 34860 6690 34916 7196
rect 34860 6638 34862 6690
rect 34914 6638 34916 6690
rect 34860 6626 34916 6638
rect 34636 5854 34638 5906
rect 34690 5854 34692 5906
rect 34636 4338 34692 5854
rect 34972 5122 35028 10332
rect 35084 8260 35140 11452
rect 35420 10834 35476 11564
rect 35420 10782 35422 10834
rect 35474 10782 35476 10834
rect 35420 10770 35476 10782
rect 35532 10612 35588 10622
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 9938 35476 9950
rect 35420 9886 35422 9938
rect 35474 9886 35476 9938
rect 35420 9716 35476 9886
rect 35420 9650 35476 9660
rect 35420 9156 35476 9166
rect 35420 9062 35476 9100
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35532 8482 35588 10556
rect 35644 9716 35700 12014
rect 35756 11732 35812 13580
rect 35868 13634 35924 13646
rect 35868 13582 35870 13634
rect 35922 13582 35924 13634
rect 35868 12516 35924 13582
rect 35868 12450 35924 12460
rect 35980 13186 36036 13198
rect 35980 13134 35982 13186
rect 36034 13134 36036 13186
rect 35980 12738 36036 13134
rect 35980 12686 35982 12738
rect 36034 12686 36036 12738
rect 35756 11666 35812 11676
rect 35980 12068 36036 12686
rect 36428 12740 36484 12750
rect 36428 12646 36484 12684
rect 36540 12402 36596 15372
rect 36540 12350 36542 12402
rect 36594 12350 36596 12402
rect 36540 12338 36596 12350
rect 36652 12740 36708 12750
rect 36092 12068 36148 12078
rect 35980 12066 36148 12068
rect 35980 12014 36094 12066
rect 36146 12014 36148 12066
rect 35980 12012 36148 12014
rect 35868 10612 35924 10622
rect 35644 9650 35700 9660
rect 35756 10610 35924 10612
rect 35756 10558 35870 10610
rect 35922 10558 35924 10610
rect 35756 10556 35924 10558
rect 35532 8430 35534 8482
rect 35586 8430 35588 8482
rect 35532 8418 35588 8430
rect 35644 9044 35700 9054
rect 35084 8194 35140 8204
rect 35644 8258 35700 8988
rect 35644 8206 35646 8258
rect 35698 8206 35700 8258
rect 35644 8194 35700 8206
rect 35532 8034 35588 8046
rect 35532 7982 35534 8034
rect 35586 7982 35588 8034
rect 35532 7924 35588 7982
rect 35532 7858 35588 7868
rect 35532 7588 35588 7598
rect 35532 7494 35588 7532
rect 35084 7252 35140 7262
rect 35084 6690 35140 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6638 35086 6690
rect 35138 6638 35140 6690
rect 35084 6626 35140 6638
rect 35532 6692 35588 6702
rect 35756 6692 35812 10556
rect 35868 10546 35924 10556
rect 35980 10164 36036 12012
rect 36092 12002 36148 12012
rect 36540 12068 36596 12078
rect 36204 11732 36260 11742
rect 36092 10836 36148 10846
rect 36092 10388 36148 10780
rect 36204 10722 36260 11676
rect 36204 10670 36206 10722
rect 36258 10670 36260 10722
rect 36204 10658 36260 10670
rect 36092 10322 36148 10332
rect 36092 10164 36148 10174
rect 35980 10108 36092 10164
rect 35532 6690 35812 6692
rect 35532 6638 35534 6690
rect 35586 6638 35812 6690
rect 35532 6636 35812 6638
rect 35868 9602 35924 9614
rect 35868 9550 35870 9602
rect 35922 9550 35924 9602
rect 35532 6626 35588 6636
rect 35308 6466 35364 6478
rect 35308 6414 35310 6466
rect 35362 6414 35364 6466
rect 35308 6020 35364 6414
rect 35420 6020 35476 6030
rect 35308 6018 35476 6020
rect 35308 5966 35422 6018
rect 35474 5966 35476 6018
rect 35308 5964 35476 5966
rect 35420 5954 35476 5964
rect 35868 6020 35924 9550
rect 36092 9602 36148 10108
rect 36092 9550 36094 9602
rect 36146 9550 36148 9602
rect 36092 9044 36148 9550
rect 36092 8978 36148 8988
rect 36204 9828 36260 9838
rect 36204 8820 36260 9772
rect 36204 8754 36260 8764
rect 36316 9716 36372 9726
rect 36092 8596 36148 8606
rect 36092 6802 36148 8540
rect 36204 8260 36260 8270
rect 36316 8260 36372 9660
rect 36204 8258 36372 8260
rect 36204 8206 36206 8258
rect 36258 8206 36372 8258
rect 36204 8204 36372 8206
rect 36540 8258 36596 12012
rect 36540 8206 36542 8258
rect 36594 8206 36596 8258
rect 36204 8194 36260 8204
rect 36540 8194 36596 8206
rect 36652 9602 36708 12684
rect 37436 12738 37492 12750
rect 37884 12740 37940 12750
rect 37436 12686 37438 12738
rect 37490 12686 37492 12738
rect 36764 12068 36820 12078
rect 36764 11506 36820 12012
rect 36988 12066 37044 12078
rect 36988 12014 36990 12066
rect 37042 12014 37044 12066
rect 36988 11732 37044 12014
rect 37436 11844 37492 12686
rect 37436 11778 37492 11788
rect 37772 12738 37940 12740
rect 37772 12686 37886 12738
rect 37938 12686 37940 12738
rect 37772 12684 37940 12686
rect 36988 11666 37044 11676
rect 37772 11732 37828 12684
rect 37884 12674 37940 12684
rect 40572 12740 40628 22094
rect 40460 12404 40516 12414
rect 40572 12404 40628 12684
rect 42140 14644 42196 14654
rect 42028 12516 42084 12526
rect 41468 12404 41524 12414
rect 40460 12402 41524 12404
rect 40460 12350 40462 12402
rect 40514 12350 41470 12402
rect 41522 12350 41524 12402
rect 40460 12348 41524 12350
rect 40460 12338 40516 12348
rect 37884 12068 37940 12078
rect 37884 11974 37940 12012
rect 37996 12068 38052 12078
rect 38556 12068 38612 12078
rect 37996 12066 38612 12068
rect 37996 12014 37998 12066
rect 38050 12014 38558 12066
rect 38610 12014 38612 12066
rect 37996 12012 38612 12014
rect 37996 12002 38052 12012
rect 36764 11454 36766 11506
rect 36818 11454 36820 11506
rect 36764 11442 36820 11454
rect 37660 11396 37716 11406
rect 37660 11302 37716 11340
rect 37548 11284 37604 11294
rect 37548 11190 37604 11228
rect 36876 10724 36932 10734
rect 36876 10630 36932 10668
rect 36988 10610 37044 10622
rect 36988 10558 36990 10610
rect 37042 10558 37044 10610
rect 36652 9550 36654 9602
rect 36706 9550 36708 9602
rect 36316 8036 36372 8046
rect 36316 7942 36372 7980
rect 36092 6750 36094 6802
rect 36146 6750 36148 6802
rect 36092 6738 36148 6750
rect 36204 7924 36260 7934
rect 35980 6692 36036 6702
rect 35980 6598 36036 6636
rect 35868 5954 35924 5964
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35980 5348 36036 5358
rect 35980 5254 36036 5292
rect 34972 5070 34974 5122
rect 35026 5070 35028 5122
rect 34972 5058 35028 5070
rect 35420 5124 35476 5134
rect 35084 5012 35140 5022
rect 35084 4918 35140 4956
rect 35420 5010 35476 5068
rect 35420 4958 35422 5010
rect 35474 4958 35476 5010
rect 35420 4946 35476 4958
rect 36092 5012 36148 5022
rect 36204 5012 36260 7868
rect 36428 7700 36484 7710
rect 36316 7252 36372 7262
rect 36316 6914 36372 7196
rect 36316 6862 36318 6914
rect 36370 6862 36372 6914
rect 36316 6850 36372 6862
rect 36316 5348 36372 5358
rect 36428 5348 36484 7644
rect 36316 5346 36484 5348
rect 36316 5294 36318 5346
rect 36370 5294 36484 5346
rect 36316 5292 36484 5294
rect 36652 6916 36708 9550
rect 36876 10386 36932 10398
rect 36876 10334 36878 10386
rect 36930 10334 36932 10386
rect 36876 7364 36932 10334
rect 36988 10164 37044 10558
rect 36988 10098 37044 10108
rect 37436 10498 37492 10510
rect 37436 10446 37438 10498
rect 37490 10446 37492 10498
rect 37436 10164 37492 10446
rect 37772 10500 37828 11676
rect 37996 11844 38052 11854
rect 37772 10434 37828 10444
rect 37884 11394 37940 11406
rect 37884 11342 37886 11394
rect 37938 11342 37940 11394
rect 37884 10388 37940 11342
rect 37996 11394 38052 11788
rect 37996 11342 37998 11394
rect 38050 11342 38052 11394
rect 37996 11060 38052 11342
rect 37996 11004 38500 11060
rect 38220 10836 38276 10846
rect 38276 10780 38388 10836
rect 38220 10742 38276 10780
rect 37996 10612 38052 10622
rect 37996 10518 38052 10556
rect 38220 10498 38276 10510
rect 38220 10446 38222 10498
rect 38274 10446 38276 10498
rect 38220 10388 38276 10446
rect 37884 10332 38276 10388
rect 37436 10098 37492 10108
rect 37660 9940 37716 9950
rect 37660 9846 37716 9884
rect 37884 9826 37940 9838
rect 37884 9774 37886 9826
rect 37938 9774 37940 9826
rect 37548 9714 37604 9726
rect 37548 9662 37550 9714
rect 37602 9662 37604 9714
rect 37436 9380 37492 9390
rect 37436 8484 37492 9324
rect 37548 9156 37604 9662
rect 37884 9380 37940 9774
rect 38108 9828 38164 9838
rect 38108 9492 38164 9772
rect 38220 9716 38276 10332
rect 38220 9650 38276 9660
rect 38108 9436 38276 9492
rect 38220 9380 38276 9436
rect 37884 9324 38164 9380
rect 37548 9090 37604 9100
rect 38108 9154 38164 9324
rect 38220 9314 38276 9324
rect 38108 9102 38110 9154
rect 38162 9102 38164 9154
rect 38108 9090 38164 9102
rect 38220 9044 38276 9054
rect 38332 9044 38388 10780
rect 38444 9828 38500 11004
rect 38556 10612 38612 12012
rect 38892 12066 38948 12078
rect 38892 12014 38894 12066
rect 38946 12014 38948 12066
rect 38892 11508 38948 12014
rect 38780 11452 38948 11508
rect 39564 12066 39620 12078
rect 39564 12014 39566 12066
rect 39618 12014 39620 12066
rect 38668 11396 38724 11406
rect 38668 11302 38724 11340
rect 38556 10546 38612 10556
rect 38780 10498 38836 11452
rect 38780 10446 38782 10498
rect 38834 10446 38836 10498
rect 38780 10052 38836 10446
rect 38780 9986 38836 9996
rect 39004 11396 39060 11406
rect 39004 10612 39060 11340
rect 39228 11394 39284 11406
rect 39228 11342 39230 11394
rect 39282 11342 39284 11394
rect 39228 10836 39284 11342
rect 39228 10770 39284 10780
rect 39564 10836 39620 12014
rect 40796 11618 40852 11630
rect 40796 11566 40798 11618
rect 40850 11566 40852 11618
rect 39676 11396 39732 11406
rect 39676 11172 39732 11340
rect 40348 11172 40404 11182
rect 40796 11172 40852 11566
rect 39676 11170 39844 11172
rect 39676 11118 39678 11170
rect 39730 11118 39844 11170
rect 39676 11116 39844 11118
rect 39676 11106 39732 11116
rect 39564 10770 39620 10780
rect 38668 9940 38724 9950
rect 39004 9940 39060 10556
rect 38668 9846 38724 9884
rect 38892 9884 39060 9940
rect 39116 10724 39172 10734
rect 38444 9762 38500 9772
rect 38780 9716 38836 9726
rect 38780 9622 38836 9660
rect 38556 9604 38612 9614
rect 38220 9042 38388 9044
rect 38220 8990 38222 9042
rect 38274 8990 38388 9042
rect 38220 8988 38388 8990
rect 38444 9044 38500 9054
rect 37548 8932 37604 8942
rect 37548 8838 37604 8876
rect 37996 8596 38052 8606
rect 37548 8484 37604 8494
rect 37436 8482 37604 8484
rect 37436 8430 37550 8482
rect 37602 8430 37604 8482
rect 37436 8428 37604 8430
rect 37548 8418 37604 8428
rect 37660 8034 37716 8046
rect 37660 7982 37662 8034
rect 37714 7982 37716 8034
rect 37660 7588 37716 7982
rect 37660 7522 37716 7532
rect 37772 8034 37828 8046
rect 37772 7982 37774 8034
rect 37826 7982 37828 8034
rect 36876 7298 36932 7308
rect 37660 7364 37716 7374
rect 37660 7270 37716 7308
rect 36316 5282 36372 5292
rect 36652 5236 36708 6860
rect 36764 6804 36820 6814
rect 36764 6710 36820 6748
rect 37772 6802 37828 7982
rect 37772 6750 37774 6802
rect 37826 6750 37828 6802
rect 37772 6738 37828 6750
rect 37884 7476 37940 7486
rect 37884 6690 37940 7420
rect 37884 6638 37886 6690
rect 37938 6638 37940 6690
rect 37884 6626 37940 6638
rect 37660 6468 37716 6478
rect 37996 6468 38052 8540
rect 38220 8484 38276 8988
rect 38444 8950 38500 8988
rect 38108 8428 38276 8484
rect 38108 6580 38164 8428
rect 38556 8146 38612 9548
rect 38892 9492 38948 9884
rect 38668 9436 38948 9492
rect 39004 9716 39060 9726
rect 38668 9042 38724 9436
rect 38668 8990 38670 9042
rect 38722 8990 38724 9042
rect 38668 8978 38724 8990
rect 39004 8932 39060 9660
rect 39116 9268 39172 10668
rect 39788 10612 39844 11116
rect 40348 11170 40852 11172
rect 40348 11118 40350 11170
rect 40402 11118 40798 11170
rect 40850 11118 40852 11170
rect 40348 11116 40852 11118
rect 40348 11106 40404 11116
rect 40236 10836 40292 10846
rect 39788 10546 39844 10556
rect 40124 10612 40180 10622
rect 40124 10518 40180 10556
rect 39228 10498 39284 10510
rect 39228 10446 39230 10498
rect 39282 10446 39284 10498
rect 39228 10276 39284 10446
rect 39676 10498 39732 10510
rect 39676 10446 39678 10498
rect 39730 10446 39732 10498
rect 39676 10388 39732 10446
rect 39676 10322 39732 10332
rect 39228 10210 39284 10220
rect 39788 10276 39844 10286
rect 39564 9716 39620 9726
rect 39564 9622 39620 9660
rect 39676 9602 39732 9614
rect 39676 9550 39678 9602
rect 39730 9550 39732 9602
rect 39228 9268 39284 9278
rect 39116 9266 39284 9268
rect 39116 9214 39230 9266
rect 39282 9214 39284 9266
rect 39116 9212 39284 9214
rect 39228 9202 39284 9212
rect 39676 9044 39732 9550
rect 39788 9266 39844 10220
rect 40124 9828 40180 9838
rect 40124 9734 40180 9772
rect 39788 9214 39790 9266
rect 39842 9214 39844 9266
rect 39788 9202 39844 9214
rect 40236 9266 40292 10780
rect 40236 9214 40238 9266
rect 40290 9214 40292 9266
rect 39676 8978 39732 8988
rect 40012 9044 40068 9054
rect 39004 8866 39060 8876
rect 39340 8930 39396 8942
rect 39340 8878 39342 8930
rect 39394 8878 39396 8930
rect 38668 8820 38724 8830
rect 38668 8258 38724 8764
rect 39340 8596 39396 8878
rect 39340 8530 39396 8540
rect 39564 8372 39620 8382
rect 39564 8278 39620 8316
rect 38668 8206 38670 8258
rect 38722 8206 38724 8258
rect 38668 8194 38724 8206
rect 39228 8260 39284 8270
rect 39228 8166 39284 8204
rect 38556 8094 38558 8146
rect 38610 8094 38612 8146
rect 38556 8082 38612 8094
rect 38220 8036 38276 8046
rect 38220 7586 38276 7980
rect 38332 8036 38388 8046
rect 38332 8034 38500 8036
rect 38332 7982 38334 8034
rect 38386 7982 38500 8034
rect 38332 7980 38500 7982
rect 38332 7970 38388 7980
rect 38332 7700 38388 7710
rect 38332 7606 38388 7644
rect 38220 7534 38222 7586
rect 38274 7534 38276 7586
rect 38220 7522 38276 7534
rect 38108 6578 38276 6580
rect 38108 6526 38110 6578
rect 38162 6526 38276 6578
rect 38108 6524 38276 6526
rect 38108 6514 38164 6524
rect 37660 6466 38052 6468
rect 37660 6414 37662 6466
rect 37714 6414 38052 6466
rect 37660 6412 38052 6414
rect 37660 6402 37716 6412
rect 37660 6132 37716 6142
rect 37548 6020 37604 6030
rect 37436 5908 37492 5918
rect 36764 5236 36820 5246
rect 36652 5234 36820 5236
rect 36652 5182 36766 5234
rect 36818 5182 36820 5234
rect 36652 5180 36820 5182
rect 37436 5236 37492 5852
rect 37548 5794 37604 5964
rect 37548 5742 37550 5794
rect 37602 5742 37604 5794
rect 37548 5730 37604 5742
rect 37548 5236 37604 5246
rect 37436 5234 37604 5236
rect 37436 5182 37550 5234
rect 37602 5182 37604 5234
rect 37436 5180 37604 5182
rect 36764 5170 36820 5180
rect 37548 5170 37604 5180
rect 36092 5010 36260 5012
rect 36092 4958 36094 5010
rect 36146 4958 36260 5010
rect 36092 4956 36260 4958
rect 36092 4946 36148 4956
rect 35308 4898 35364 4910
rect 35308 4846 35310 4898
rect 35362 4846 35364 4898
rect 35308 4452 35364 4846
rect 35420 4452 35476 4462
rect 35308 4450 35476 4452
rect 35308 4398 35422 4450
rect 35474 4398 35476 4450
rect 35308 4396 35476 4398
rect 35420 4386 35476 4396
rect 34636 4286 34638 4338
rect 34690 4286 34692 4338
rect 34636 4274 34692 4286
rect 36092 4228 36148 4238
rect 34524 4060 35028 4116
rect 33852 3668 33908 3678
rect 33852 3574 33908 3612
rect 33180 3556 33236 3566
rect 33068 3554 33236 3556
rect 33068 3502 33182 3554
rect 33234 3502 33236 3554
rect 33068 3500 33236 3502
rect 33180 3490 33236 3500
rect 33404 3556 33460 3566
rect 32060 1708 32228 1764
rect 32060 800 32116 1708
rect 33404 800 33460 3500
rect 34972 3554 35028 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34972 3502 34974 3554
rect 35026 3502 35028 3554
rect 34972 3490 35028 3502
rect 35644 3666 35700 3678
rect 35644 3614 35646 3666
rect 35698 3614 35700 3666
rect 35644 3556 35700 3614
rect 35644 3490 35700 3500
rect 34748 3444 34804 3454
rect 34748 800 34804 3388
rect 36092 800 36148 4172
rect 37548 4228 37604 4238
rect 37660 4228 37716 6076
rect 38108 6132 38164 6142
rect 38108 5906 38164 6076
rect 38220 6130 38276 6524
rect 38220 6078 38222 6130
rect 38274 6078 38276 6130
rect 38220 6066 38276 6078
rect 38108 5854 38110 5906
rect 38162 5854 38164 5906
rect 38108 5842 38164 5854
rect 38332 5684 38388 5694
rect 37884 5348 37940 5358
rect 37884 5234 37940 5292
rect 37884 5182 37886 5234
rect 37938 5182 37940 5234
rect 37884 5124 37940 5182
rect 38332 5234 38388 5628
rect 38444 5348 38500 7980
rect 39452 8034 39508 8046
rect 39452 7982 39454 8034
rect 39506 7982 39508 8034
rect 38556 7476 38612 7486
rect 38556 5962 38612 7420
rect 39228 7362 39284 7374
rect 39228 7310 39230 7362
rect 39282 7310 39284 7362
rect 39004 6580 39060 6590
rect 39004 6578 39172 6580
rect 39004 6526 39006 6578
rect 39058 6526 39172 6578
rect 39004 6524 39172 6526
rect 39004 6514 39060 6524
rect 38556 5910 38558 5962
rect 38610 5910 38612 5962
rect 38556 5898 38612 5910
rect 38444 5282 38500 5292
rect 38332 5182 38334 5234
rect 38386 5182 38388 5234
rect 38332 5170 38388 5182
rect 37884 5058 37940 5068
rect 39004 5012 39060 5022
rect 38780 5010 39060 5012
rect 38780 4958 39006 5010
rect 39058 4958 39060 5010
rect 38780 4956 39060 4958
rect 37548 4226 37716 4228
rect 37548 4174 37550 4226
rect 37602 4174 37716 4226
rect 37548 4172 37716 4174
rect 38220 4228 38276 4238
rect 37548 4162 37604 4172
rect 38220 4134 38276 4172
rect 38332 4116 38388 4126
rect 38332 3554 38388 4060
rect 38332 3502 38334 3554
rect 38386 3502 38388 3554
rect 38332 3490 38388 3502
rect 37212 3444 37268 3482
rect 37212 3378 37268 3388
rect 37436 3444 37492 3454
rect 37436 800 37492 3388
rect 38780 800 38836 4956
rect 39004 4946 39060 4956
rect 39116 3668 39172 6524
rect 39228 3892 39284 7310
rect 39340 5908 39396 5918
rect 39340 5814 39396 5852
rect 39452 5124 39508 7982
rect 39788 7924 39844 7934
rect 39788 7588 39844 7868
rect 39676 7364 39732 7374
rect 39564 6020 39620 6030
rect 39564 5926 39620 5964
rect 39676 5684 39732 7308
rect 39788 5796 39844 7532
rect 40012 6020 40068 8988
rect 40124 8372 40180 8382
rect 40236 8372 40292 9214
rect 40460 8484 40516 11116
rect 40796 11106 40852 11116
rect 41244 11172 41300 11182
rect 41244 11170 41412 11172
rect 41244 11118 41246 11170
rect 41298 11118 41412 11170
rect 41244 11116 41412 11118
rect 41244 11106 41300 11116
rect 40572 10836 40628 10846
rect 40572 10742 40628 10780
rect 41356 10612 41412 11116
rect 40572 10052 40628 10062
rect 40572 9938 40628 9996
rect 40572 9886 40574 9938
rect 40626 9886 40628 9938
rect 40572 9874 40628 9886
rect 41020 9828 41076 9838
rect 41020 9734 41076 9772
rect 40684 8930 40740 8942
rect 40684 8878 40686 8930
rect 40738 8878 40740 8930
rect 40684 8484 40740 8878
rect 40460 8372 40628 8428
rect 40684 8418 40740 8428
rect 40236 8316 40404 8372
rect 40124 8278 40180 8316
rect 40236 8146 40292 8158
rect 40236 8094 40238 8146
rect 40290 8094 40292 8146
rect 40236 7700 40292 8094
rect 40348 7924 40404 8316
rect 40572 8260 40628 8372
rect 41244 8372 41300 8382
rect 40572 8204 40964 8260
rect 40684 8036 40740 8046
rect 40684 7942 40740 7980
rect 40348 7858 40404 7868
rect 40236 7634 40292 7644
rect 40124 7476 40180 7486
rect 40124 7474 40292 7476
rect 40124 7422 40126 7474
rect 40178 7422 40292 7474
rect 40124 7420 40292 7422
rect 40124 7410 40180 7420
rect 40124 6692 40180 6702
rect 40124 6598 40180 6636
rect 40236 6130 40292 7420
rect 40684 7364 40740 7374
rect 40236 6078 40238 6130
rect 40290 6078 40292 6130
rect 40236 6066 40292 6078
rect 40348 7362 40740 7364
rect 40348 7310 40686 7362
rect 40738 7310 40740 7362
rect 40348 7308 40740 7310
rect 40124 6020 40180 6030
rect 40012 6018 40180 6020
rect 40012 5966 40126 6018
rect 40178 5966 40180 6018
rect 40012 5964 40180 5966
rect 40124 5954 40180 5964
rect 40348 6020 40404 7308
rect 40684 7298 40740 7308
rect 40796 7252 40852 7262
rect 40796 7158 40852 7196
rect 40796 6692 40852 6702
rect 40908 6692 40964 8204
rect 41132 8148 41188 8158
rect 41132 8054 41188 8092
rect 40348 5954 40404 5964
rect 40460 6690 40964 6692
rect 40460 6638 40798 6690
rect 40850 6638 40964 6690
rect 40460 6636 40964 6638
rect 40460 5906 40516 6636
rect 40796 6626 40852 6636
rect 40908 6132 40964 6636
rect 40908 6066 40964 6076
rect 41020 8036 41076 8046
rect 41020 6804 41076 7980
rect 40460 5854 40462 5906
rect 40514 5854 40516 5906
rect 40460 5842 40516 5854
rect 39788 5740 40292 5796
rect 39676 5628 39956 5684
rect 39452 5058 39508 5068
rect 39900 5122 39956 5628
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 5058 39956 5070
rect 40124 5236 40180 5246
rect 40012 4564 40068 4574
rect 40012 4470 40068 4508
rect 39340 4452 39396 4462
rect 39340 4338 39396 4396
rect 39340 4286 39342 4338
rect 39394 4286 39396 4338
rect 39340 4274 39396 4286
rect 39900 4116 39956 4126
rect 39900 4022 39956 4060
rect 39228 3826 39284 3836
rect 40124 3780 40180 5180
rect 40236 4450 40292 5740
rect 40684 5124 40740 5134
rect 40684 5030 40740 5068
rect 41020 4900 41076 6748
rect 40684 4844 41076 4900
rect 41244 6802 41300 8316
rect 41244 6750 41246 6802
rect 41298 6750 41300 6802
rect 40684 4562 40740 4844
rect 40684 4510 40686 4562
rect 40738 4510 40740 4562
rect 40684 4498 40740 4510
rect 41244 4564 41300 6750
rect 41356 6468 41412 10556
rect 41468 10834 41524 12348
rect 42028 12402 42084 12460
rect 42028 12350 42030 12402
rect 42082 12350 42084 12402
rect 42028 12338 42084 12350
rect 41692 11618 41748 11630
rect 41692 11566 41694 11618
rect 41746 11566 41748 11618
rect 41692 11506 41748 11566
rect 41692 11454 41694 11506
rect 41746 11454 41748 11506
rect 41692 11442 41748 11454
rect 41468 10782 41470 10834
rect 41522 10782 41524 10834
rect 41468 9938 41524 10782
rect 41804 10500 41860 10510
rect 41916 10500 41972 10510
rect 41860 10498 41972 10500
rect 41860 10446 41918 10498
rect 41970 10446 41972 10498
rect 41860 10444 41972 10446
rect 41468 9886 41470 9938
rect 41522 9886 41524 9938
rect 41468 9266 41524 9886
rect 41468 9214 41470 9266
rect 41522 9214 41524 9266
rect 41468 8372 41524 9214
rect 41468 7812 41524 8316
rect 41580 10164 41636 10174
rect 41580 8370 41636 10108
rect 41804 8428 41860 10444
rect 41916 10434 41972 10444
rect 41916 10276 41972 10286
rect 41916 9938 41972 10220
rect 41916 9886 41918 9938
rect 41970 9886 41972 9938
rect 41916 9874 41972 9886
rect 41916 9604 41972 9614
rect 41916 9266 41972 9548
rect 41916 9214 41918 9266
rect 41970 9214 41972 9266
rect 41916 9202 41972 9214
rect 41804 8372 41972 8428
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 41468 7756 41860 7812
rect 41804 7698 41860 7756
rect 41804 7646 41806 7698
rect 41858 7646 41860 7698
rect 41804 7634 41860 7646
rect 41692 7364 41748 7374
rect 41692 7270 41748 7308
rect 41580 7252 41636 7262
rect 41580 7158 41636 7196
rect 41692 6692 41748 6702
rect 41356 6412 41636 6468
rect 41580 6018 41636 6412
rect 41692 6130 41748 6636
rect 41916 6690 41972 8372
rect 42028 8036 42084 8046
rect 42028 7942 42084 7980
rect 41916 6638 41918 6690
rect 41970 6638 41972 6690
rect 41916 6244 41972 6638
rect 41916 6178 41972 6188
rect 42028 6468 42084 6478
rect 41692 6078 41694 6130
rect 41746 6078 41748 6130
rect 41692 6066 41748 6078
rect 41804 6132 41860 6142
rect 41804 6038 41860 6076
rect 41580 5966 41582 6018
rect 41634 5966 41636 6018
rect 41580 5954 41636 5966
rect 41804 5348 41860 5358
rect 41356 5236 41412 5246
rect 41356 5142 41412 5180
rect 41244 4498 41300 4508
rect 41692 4564 41748 4574
rect 40236 4398 40238 4450
rect 40290 4398 40292 4450
rect 40236 4386 40292 4398
rect 41580 4452 41636 4462
rect 41580 4358 41636 4396
rect 39116 3602 39172 3612
rect 40012 3724 40180 3780
rect 40908 3780 40964 3790
rect 39004 3444 39060 3454
rect 39004 3350 39060 3388
rect 40012 2548 40068 3724
rect 40908 3666 40964 3724
rect 40908 3614 40910 3666
rect 40962 3614 40964 3666
rect 40908 3602 40964 3614
rect 41468 3668 41524 3678
rect 40124 3556 40180 3566
rect 40124 3462 40180 3500
rect 40012 2492 40180 2548
rect 40124 800 40180 2492
rect 41468 800 41524 3612
rect 41580 3666 41636 3678
rect 41580 3614 41582 3666
rect 41634 3614 41636 3666
rect 41580 3556 41636 3614
rect 41580 3490 41636 3500
rect 41692 3442 41748 4508
rect 41804 4338 41860 5292
rect 41804 4286 41806 4338
rect 41858 4286 41860 4338
rect 41804 4274 41860 4286
rect 41916 5012 41972 5022
rect 42028 5012 42084 6412
rect 41972 4956 42084 5012
rect 41916 3778 41972 4956
rect 42140 4676 42196 14588
rect 42252 6580 42308 22428
rect 42476 19908 42532 19918
rect 42364 19796 42420 19806
rect 42364 6804 42420 19740
rect 42364 6738 42420 6748
rect 42252 6524 42420 6580
rect 42140 4610 42196 4620
rect 41916 3726 41918 3778
rect 41970 3726 41972 3778
rect 41916 3714 41972 3726
rect 41692 3390 41694 3442
rect 41746 3390 41748 3442
rect 41692 3378 41748 3390
rect 42364 2996 42420 6524
rect 42364 2930 42420 2940
rect 42476 2884 42532 19852
rect 42588 3332 42644 22540
rect 42588 3266 42644 3276
rect 42476 2818 42532 2828
rect 42700 2660 42756 23884
rect 42812 12516 42868 12526
rect 42812 6468 42868 12460
rect 42812 6402 42868 6412
rect 42924 6804 42980 6814
rect 42700 2594 42756 2604
rect 42812 3892 42868 3902
rect 42812 800 42868 3836
rect 42924 2548 42980 6748
rect 42924 2482 42980 2492
rect 18844 700 19348 756
rect 19936 0 20048 800
rect 21280 0 21392 800
rect 22624 0 22736 800
rect 23968 0 24080 800
rect 25312 0 25424 800
rect 26656 0 26768 800
rect 28000 0 28112 800
rect 29344 0 29456 800
rect 30688 0 30800 800
rect 32032 0 32144 800
rect 33376 0 33488 800
rect 34720 0 34832 800
rect 36064 0 36176 800
rect 37408 0 37520 800
rect 38752 0 38864 800
rect 40096 0 40208 800
rect 41440 0 41552 800
rect 42784 0 42896 800
<< via2 >>
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 15932 32284 15988 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 2492 25506 2548 25508
rect 2492 25454 2494 25506
rect 2494 25454 2546 25506
rect 2546 25454 2548 25506
rect 2492 25452 2548 25454
rect 1708 25340 1764 25396
rect 1484 25228 1540 25284
rect 1372 23660 1428 23716
rect 1148 23548 1204 23604
rect 1036 16716 1092 16772
rect 1148 11340 1204 11396
rect 1260 22316 1316 22372
rect 1260 5964 1316 6020
rect 1484 6524 1540 6580
rect 1596 23772 1652 23828
rect 1372 5068 1428 5124
rect 13468 25340 13524 25396
rect 2940 25282 2996 25284
rect 2940 25230 2942 25282
rect 2942 25230 2994 25282
rect 2994 25230 2996 25282
rect 2940 25228 2996 25230
rect 2268 24722 2324 24724
rect 2268 24670 2270 24722
rect 2270 24670 2322 24722
rect 2322 24670 2324 24722
rect 2268 24668 2324 24670
rect 1932 23714 1988 23716
rect 1932 23662 1934 23714
rect 1934 23662 1986 23714
rect 1986 23662 1988 23714
rect 1932 23660 1988 23662
rect 2156 23378 2212 23380
rect 2156 23326 2158 23378
rect 2158 23326 2210 23378
rect 2210 23326 2212 23378
rect 2156 23324 2212 23326
rect 1820 23042 1876 23044
rect 1820 22990 1822 23042
rect 1822 22990 1874 23042
rect 1874 22990 1876 23042
rect 1820 22988 1876 22990
rect 1820 22540 1876 22596
rect 2716 24610 2772 24612
rect 2716 24558 2718 24610
rect 2718 24558 2770 24610
rect 2770 24558 2772 24610
rect 2716 24556 2772 24558
rect 3276 23884 3332 23940
rect 3836 24444 3892 24500
rect 3724 23826 3780 23828
rect 3724 23774 3726 23826
rect 3726 23774 3778 23826
rect 3778 23774 3780 23826
rect 3724 23772 3780 23774
rect 2156 22146 2212 22148
rect 2156 22094 2158 22146
rect 2158 22094 2210 22146
rect 2210 22094 2212 22146
rect 2156 22092 2212 22094
rect 2044 20690 2100 20692
rect 2044 20638 2046 20690
rect 2046 20638 2098 20690
rect 2098 20638 2100 20690
rect 2044 20636 2100 20638
rect 1932 19404 1988 19460
rect 1708 18284 1764 18340
rect 1820 18450 1876 18452
rect 1820 18398 1822 18450
rect 1822 18398 1874 18450
rect 1874 18398 1876 18450
rect 1820 18396 1876 18398
rect 2716 23100 2772 23156
rect 2604 23042 2660 23044
rect 2604 22990 2606 23042
rect 2606 22990 2658 23042
rect 2658 22990 2660 23042
rect 2604 22988 2660 22990
rect 3276 23548 3332 23604
rect 3052 23324 3108 23380
rect 3164 22876 3220 22932
rect 2380 20188 2436 20244
rect 2716 20242 2772 20244
rect 2716 20190 2718 20242
rect 2718 20190 2770 20242
rect 2770 20190 2772 20242
rect 2716 20188 2772 20190
rect 2492 19964 2548 20020
rect 2268 19122 2324 19124
rect 2268 19070 2270 19122
rect 2270 19070 2322 19122
rect 2322 19070 2324 19122
rect 2268 19068 2324 19070
rect 2828 19964 2884 20020
rect 2940 20524 2996 20580
rect 2492 19068 2548 19124
rect 2156 18956 2212 19012
rect 2156 18338 2212 18340
rect 2156 18286 2158 18338
rect 2158 18286 2210 18338
rect 2210 18286 2212 18338
rect 2156 18284 2212 18286
rect 2380 18172 2436 18228
rect 2044 17106 2100 17108
rect 2044 17054 2046 17106
rect 2046 17054 2098 17106
rect 2098 17054 2100 17106
rect 2044 17052 2100 17054
rect 1932 16994 1988 16996
rect 1932 16942 1934 16994
rect 1934 16942 1986 16994
rect 1986 16942 1988 16994
rect 1932 16940 1988 16942
rect 1708 16828 1764 16884
rect 1820 16098 1876 16100
rect 1820 16046 1822 16098
rect 1822 16046 1874 16098
rect 1874 16046 1876 16098
rect 1820 16044 1876 16046
rect 2268 16604 2324 16660
rect 2716 19010 2772 19012
rect 2716 18958 2718 19010
rect 2718 18958 2770 19010
rect 2770 18958 2772 19010
rect 2716 18956 2772 18958
rect 2716 17724 2772 17780
rect 2604 17666 2660 17668
rect 2604 17614 2606 17666
rect 2606 17614 2658 17666
rect 2658 17614 2660 17666
rect 2604 17612 2660 17614
rect 2828 17500 2884 17556
rect 1932 15260 1988 15316
rect 2268 15820 2324 15876
rect 2380 15708 2436 15764
rect 2156 14642 2212 14644
rect 2156 14590 2158 14642
rect 2158 14590 2210 14642
rect 2210 14590 2212 14642
rect 2156 14588 2212 14590
rect 1932 13634 1988 13636
rect 1932 13582 1934 13634
rect 1934 13582 1986 13634
rect 1986 13582 1988 13634
rect 1932 13580 1988 13582
rect 2044 13468 2100 13524
rect 1932 12460 1988 12516
rect 1820 11676 1876 11732
rect 1932 11004 1988 11060
rect 2604 17052 2660 17108
rect 3500 21474 3556 21476
rect 3500 21422 3502 21474
rect 3502 21422 3554 21474
rect 3554 21422 3556 21474
rect 3500 21420 3556 21422
rect 3500 20636 3556 20692
rect 3276 20188 3332 20244
rect 3164 18338 3220 18340
rect 3164 18286 3166 18338
rect 3166 18286 3218 18338
rect 3218 18286 3220 18338
rect 3164 18284 3220 18286
rect 3052 17836 3108 17892
rect 3052 17442 3108 17444
rect 3052 17390 3054 17442
rect 3054 17390 3106 17442
rect 3106 17390 3108 17442
rect 3052 17388 3108 17390
rect 2716 16994 2772 16996
rect 2716 16942 2718 16994
rect 2718 16942 2770 16994
rect 2770 16942 2772 16994
rect 2716 16940 2772 16942
rect 2828 15820 2884 15876
rect 2268 14140 2324 14196
rect 2268 12850 2324 12852
rect 2268 12798 2270 12850
rect 2270 12798 2322 12850
rect 2322 12798 2324 12850
rect 2268 12796 2324 12798
rect 2156 12236 2212 12292
rect 2492 12796 2548 12852
rect 2604 12402 2660 12404
rect 2604 12350 2606 12402
rect 2606 12350 2658 12402
rect 2658 12350 2660 12402
rect 2604 12348 2660 12350
rect 2492 11900 2548 11956
rect 2604 12124 2660 12180
rect 2380 10108 2436 10164
rect 2156 9938 2212 9940
rect 2156 9886 2158 9938
rect 2158 9886 2210 9938
rect 2210 9886 2212 9938
rect 2156 9884 2212 9886
rect 1820 9714 1876 9716
rect 1820 9662 1822 9714
rect 1822 9662 1874 9714
rect 1874 9662 1876 9714
rect 1820 9660 1876 9662
rect 3164 17052 3220 17108
rect 4956 24556 5012 24612
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4620 23714 4676 23716
rect 4620 23662 4622 23714
rect 4622 23662 4674 23714
rect 4674 23662 4676 23714
rect 4620 23660 4676 23662
rect 4396 23436 4452 23492
rect 4956 23714 5012 23716
rect 4956 23662 4958 23714
rect 4958 23662 5010 23714
rect 5010 23662 5012 23714
rect 4956 23660 5012 23662
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4844 22482 4900 22484
rect 4844 22430 4846 22482
rect 4846 22430 4898 22482
rect 4898 22430 4900 22482
rect 4844 22428 4900 22430
rect 4060 22316 4116 22372
rect 3836 21756 3892 21812
rect 4060 21756 4116 21812
rect 3836 21586 3892 21588
rect 3836 21534 3838 21586
rect 3838 21534 3890 21586
rect 3890 21534 3892 21586
rect 3836 21532 3892 21534
rect 3948 20636 4004 20692
rect 3948 20412 4004 20468
rect 3724 20300 3780 20356
rect 4732 21810 4788 21812
rect 4732 21758 4734 21810
rect 4734 21758 4786 21810
rect 4786 21758 4788 21810
rect 4732 21756 4788 21758
rect 4284 21698 4340 21700
rect 4284 21646 4286 21698
rect 4286 21646 4338 21698
rect 4338 21646 4340 21698
rect 4284 21644 4340 21646
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4732 20748 4788 20804
rect 4620 20578 4676 20580
rect 4620 20526 4622 20578
rect 4622 20526 4674 20578
rect 4674 20526 4676 20578
rect 4620 20524 4676 20526
rect 4060 20188 4116 20244
rect 3500 19404 3556 19460
rect 3388 18396 3444 18452
rect 3500 17276 3556 17332
rect 3612 19010 3668 19012
rect 3612 18958 3614 19010
rect 3614 18958 3666 19010
rect 3666 18958 3668 19010
rect 3612 18956 3668 18958
rect 4284 20188 4340 20244
rect 4060 19740 4116 19796
rect 3500 16156 3556 16212
rect 3164 15874 3220 15876
rect 3164 15822 3166 15874
rect 3166 15822 3218 15874
rect 3218 15822 3220 15874
rect 3164 15820 3220 15822
rect 3052 15538 3108 15540
rect 3052 15486 3054 15538
rect 3054 15486 3106 15538
rect 3106 15486 3108 15538
rect 3052 15484 3108 15486
rect 3052 13132 3108 13188
rect 2940 12908 2996 12964
rect 3388 15874 3444 15876
rect 3388 15822 3390 15874
rect 3390 15822 3442 15874
rect 3442 15822 3444 15874
rect 3388 15820 3444 15822
rect 3948 18060 4004 18116
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4620 18844 4676 18900
rect 4956 20860 5012 20916
rect 5068 19852 5124 19908
rect 5964 23884 6020 23940
rect 5740 23826 5796 23828
rect 5740 23774 5742 23826
rect 5742 23774 5794 23826
rect 5794 23774 5796 23826
rect 5740 23772 5796 23774
rect 5740 23324 5796 23380
rect 5404 22988 5460 23044
rect 5740 22204 5796 22260
rect 5516 22092 5572 22148
rect 5404 21586 5460 21588
rect 5404 21534 5406 21586
rect 5406 21534 5458 21586
rect 5458 21534 5460 21586
rect 5404 21532 5460 21534
rect 5740 21810 5796 21812
rect 5740 21758 5742 21810
rect 5742 21758 5794 21810
rect 5794 21758 5796 21810
rect 5740 21756 5796 21758
rect 5516 20748 5572 20804
rect 5628 21420 5684 21476
rect 6860 24722 6916 24724
rect 6860 24670 6862 24722
rect 6862 24670 6914 24722
rect 6914 24670 6916 24722
rect 6860 24668 6916 24670
rect 6412 24108 6468 24164
rect 6188 23996 6244 24052
rect 6860 23548 6916 23604
rect 6300 23100 6356 23156
rect 6860 23100 6916 23156
rect 6188 22652 6244 22708
rect 6412 22988 6468 23044
rect 6076 22428 6132 22484
rect 6300 22204 6356 22260
rect 5964 20412 6020 20468
rect 6076 20188 6132 20244
rect 5628 20076 5684 20132
rect 6300 20578 6356 20580
rect 6300 20526 6302 20578
rect 6302 20526 6354 20578
rect 6354 20526 6356 20578
rect 6300 20524 6356 20526
rect 6524 22876 6580 22932
rect 6524 21868 6580 21924
rect 6860 21868 6916 21924
rect 6412 19852 6468 19908
rect 6524 21308 6580 21364
rect 5964 19628 6020 19684
rect 5180 19404 5236 19460
rect 4284 18284 4340 18340
rect 4956 18508 5012 18564
rect 5068 18732 5124 18788
rect 4844 18284 4900 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5292 18338 5348 18340
rect 5292 18286 5294 18338
rect 5294 18286 5346 18338
rect 5346 18286 5348 18338
rect 5292 18284 5348 18286
rect 3724 16994 3780 16996
rect 3724 16942 3726 16994
rect 3726 16942 3778 16994
rect 3778 16942 3780 16994
rect 3724 16940 3780 16942
rect 3836 16882 3892 16884
rect 3836 16830 3838 16882
rect 3838 16830 3890 16882
rect 3890 16830 3892 16882
rect 3836 16828 3892 16830
rect 3948 16268 4004 16324
rect 4396 17612 4452 17668
rect 4396 17164 4452 17220
rect 5628 17666 5684 17668
rect 5628 17614 5630 17666
rect 5630 17614 5682 17666
rect 5682 17614 5684 17666
rect 5628 17612 5684 17614
rect 4844 17442 4900 17444
rect 4844 17390 4846 17442
rect 4846 17390 4898 17442
rect 4898 17390 4900 17442
rect 4844 17388 4900 17390
rect 4956 17052 5012 17108
rect 5292 17388 5348 17444
rect 5404 17276 5460 17332
rect 5068 16994 5124 16996
rect 5068 16942 5070 16994
rect 5070 16942 5122 16994
rect 5122 16942 5124 16994
rect 5068 16940 5124 16942
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16380 4900 16436
rect 3836 15820 3892 15876
rect 3612 15708 3668 15764
rect 4060 15708 4116 15764
rect 3500 14418 3556 14420
rect 3500 14366 3502 14418
rect 3502 14366 3554 14418
rect 3554 14366 3556 14418
rect 3500 14364 3556 14366
rect 3612 14306 3668 14308
rect 3612 14254 3614 14306
rect 3614 14254 3666 14306
rect 3666 14254 3668 14306
rect 3612 14252 3668 14254
rect 3276 12796 3332 12852
rect 2828 12178 2884 12180
rect 2828 12126 2830 12178
rect 2830 12126 2882 12178
rect 2882 12126 2884 12178
rect 2828 12124 2884 12126
rect 2156 9660 2212 9716
rect 1932 8482 1988 8484
rect 1932 8430 1934 8482
rect 1934 8430 1986 8482
rect 1986 8430 1988 8482
rect 1932 8428 1988 8430
rect 2044 8204 2100 8260
rect 2156 8540 2212 8596
rect 1596 4844 1652 4900
rect 1708 7980 1764 8036
rect 2268 8092 2324 8148
rect 2044 7532 2100 7588
rect 1932 7420 1988 7476
rect 1820 5234 1876 5236
rect 1820 5182 1822 5234
rect 1822 5182 1874 5234
rect 1874 5182 1876 5234
rect 1820 5180 1876 5182
rect 2716 9938 2772 9940
rect 2716 9886 2718 9938
rect 2718 9886 2770 9938
rect 2770 9886 2772 9938
rect 2716 9884 2772 9886
rect 3164 12124 3220 12180
rect 3388 12908 3444 12964
rect 3500 11900 3556 11956
rect 3276 11676 3332 11732
rect 3388 11452 3444 11508
rect 3164 11228 3220 11284
rect 3052 9772 3108 9828
rect 2940 8428 2996 8484
rect 3052 8370 3108 8372
rect 3052 8318 3054 8370
rect 3054 8318 3106 8370
rect 3106 8318 3108 8370
rect 3052 8316 3108 8318
rect 2380 7980 2436 8036
rect 3948 15148 4004 15204
rect 3836 14700 3892 14756
rect 4172 15372 4228 15428
rect 4732 16268 4788 16324
rect 4620 15820 4676 15876
rect 4508 15708 4564 15764
rect 4620 15314 4676 15316
rect 4620 15262 4622 15314
rect 4622 15262 4674 15314
rect 4674 15262 4676 15314
rect 4620 15260 4676 15262
rect 4844 15036 4900 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4396 14306 4452 14308
rect 4396 14254 4398 14306
rect 4398 14254 4450 14306
rect 4450 14254 4452 14306
rect 4396 14252 4452 14254
rect 4284 14140 4340 14196
rect 3836 13244 3892 13300
rect 3724 13020 3780 13076
rect 6748 21084 6804 21140
rect 6636 20748 6692 20804
rect 7196 21980 7252 22036
rect 7084 20914 7140 20916
rect 7084 20862 7086 20914
rect 7086 20862 7138 20914
rect 7138 20862 7140 20914
rect 7084 20860 7140 20862
rect 6636 19180 6692 19236
rect 6524 18732 6580 18788
rect 6636 18620 6692 18676
rect 6412 18562 6468 18564
rect 6412 18510 6414 18562
rect 6414 18510 6466 18562
rect 6466 18510 6468 18562
rect 6412 18508 6468 18510
rect 5964 18396 6020 18452
rect 6524 18396 6580 18452
rect 6412 18284 6468 18340
rect 5852 17948 5908 18004
rect 6300 17890 6356 17892
rect 6300 17838 6302 17890
rect 6302 17838 6354 17890
rect 6354 17838 6356 17890
rect 6300 17836 6356 17838
rect 6076 17500 6132 17556
rect 5852 17388 5908 17444
rect 5068 15932 5124 15988
rect 5516 15932 5572 15988
rect 5180 15820 5236 15876
rect 5404 15538 5460 15540
rect 5404 15486 5406 15538
rect 5406 15486 5458 15538
rect 5458 15486 5460 15538
rect 5404 15484 5460 15486
rect 4956 13916 5012 13972
rect 5404 14700 5460 14756
rect 4844 13746 4900 13748
rect 4844 13694 4846 13746
rect 4846 13694 4898 13746
rect 4898 13694 4900 13746
rect 4844 13692 4900 13694
rect 4060 13634 4116 13636
rect 4060 13582 4062 13634
rect 4062 13582 4114 13634
rect 4114 13582 4116 13634
rect 5180 13692 5236 13748
rect 4060 13580 4116 13582
rect 4844 13468 4900 13524
rect 4476 13354 4532 13356
rect 4060 13244 4116 13300
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3724 12572 3780 12628
rect 3948 12684 4004 12740
rect 3836 12348 3892 12404
rect 3948 12290 4004 12292
rect 3948 12238 3950 12290
rect 3950 12238 4002 12290
rect 4002 12238 4004 12290
rect 3948 12236 4004 12238
rect 4172 12236 4228 12292
rect 4396 12796 4452 12852
rect 3724 12178 3780 12180
rect 3724 12126 3726 12178
rect 3726 12126 3778 12178
rect 3778 12126 3780 12178
rect 3724 12124 3780 12126
rect 3612 10556 3668 10612
rect 3724 11788 3780 11844
rect 4284 12012 4340 12068
rect 5740 16322 5796 16324
rect 5740 16270 5742 16322
rect 5742 16270 5794 16322
rect 5794 16270 5796 16322
rect 5740 16268 5796 16270
rect 6636 18060 6692 18116
rect 5964 16828 6020 16884
rect 6524 16994 6580 16996
rect 6524 16942 6526 16994
rect 6526 16942 6578 16994
rect 6578 16942 6580 16994
rect 6524 16940 6580 16942
rect 6412 16716 6468 16772
rect 6076 16322 6132 16324
rect 6076 16270 6078 16322
rect 6078 16270 6130 16322
rect 6130 16270 6132 16322
rect 6076 16268 6132 16270
rect 5852 15426 5908 15428
rect 5852 15374 5854 15426
rect 5854 15374 5906 15426
rect 5906 15374 5908 15426
rect 5852 15372 5908 15374
rect 6300 15426 6356 15428
rect 6300 15374 6302 15426
rect 6302 15374 6354 15426
rect 6354 15374 6356 15426
rect 6300 15372 6356 15374
rect 6076 14924 6132 14980
rect 5740 14700 5796 14756
rect 5852 14306 5908 14308
rect 5852 14254 5854 14306
rect 5854 14254 5906 14306
rect 5906 14254 5908 14306
rect 5852 14252 5908 14254
rect 5628 13692 5684 13748
rect 4844 12908 4900 12964
rect 4732 12236 4788 12292
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4844 11676 4900 11732
rect 4396 10892 4452 10948
rect 4508 10834 4564 10836
rect 4508 10782 4510 10834
rect 4510 10782 4562 10834
rect 4562 10782 4564 10834
rect 4508 10780 4564 10782
rect 3612 10220 3668 10276
rect 3276 9996 3332 10052
rect 5404 12908 5460 12964
rect 5068 12572 5124 12628
rect 5180 12348 5236 12404
rect 4172 10556 4228 10612
rect 3948 10220 4004 10276
rect 4060 10332 4116 10388
rect 4172 9884 4228 9940
rect 3276 9212 3332 9268
rect 4172 9436 4228 9492
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4732 9884 4788 9940
rect 5180 11116 5236 11172
rect 5292 10386 5348 10388
rect 5292 10334 5294 10386
rect 5294 10334 5346 10386
rect 5346 10334 5348 10386
rect 5292 10332 5348 10334
rect 4956 10050 5012 10052
rect 4956 9998 4958 10050
rect 4958 9998 5010 10050
rect 5010 9998 5012 10050
rect 4956 9996 5012 9998
rect 4732 9324 4788 9380
rect 4284 8988 4340 9044
rect 3948 8764 4004 8820
rect 3500 8146 3556 8148
rect 3500 8094 3502 8146
rect 3502 8094 3554 8146
rect 3554 8094 3556 8146
rect 3500 8092 3556 8094
rect 2828 7756 2884 7812
rect 3724 8034 3780 8036
rect 3724 7982 3726 8034
rect 3726 7982 3778 8034
rect 3778 7982 3780 8034
rect 3724 7980 3780 7982
rect 2828 6578 2884 6580
rect 2828 6526 2830 6578
rect 2830 6526 2882 6578
rect 2882 6526 2884 6578
rect 2828 6524 2884 6526
rect 2716 6412 2772 6468
rect 2492 5010 2548 5012
rect 2492 4958 2494 5010
rect 2494 4958 2546 5010
rect 2546 4958 2548 5010
rect 2492 4956 2548 4958
rect 2156 4508 2212 4564
rect 1036 3052 1092 3108
rect 1148 2492 1204 2548
rect 2828 3164 2884 3220
rect 3500 7868 3556 7924
rect 3276 6748 3332 6804
rect 4060 8034 4116 8036
rect 4060 7982 4062 8034
rect 4062 7982 4114 8034
rect 4114 7982 4116 8034
rect 4060 7980 4116 7982
rect 4172 7308 4228 7364
rect 3500 5180 3556 5236
rect 4172 6188 4228 6244
rect 3276 4956 3332 5012
rect 3276 3724 3332 3780
rect 2268 2492 2324 2548
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4844 7868 4900 7924
rect 5404 9660 5460 9716
rect 5180 8876 5236 8932
rect 5292 8652 5348 8708
rect 5068 8146 5124 8148
rect 5068 8094 5070 8146
rect 5070 8094 5122 8146
rect 5122 8094 5124 8146
rect 5068 8092 5124 8094
rect 5740 11954 5796 11956
rect 5740 11902 5742 11954
rect 5742 11902 5794 11954
rect 5794 11902 5796 11954
rect 5740 11900 5796 11902
rect 6076 14252 6132 14308
rect 6524 15260 6580 15316
rect 6748 17052 6804 17108
rect 6860 19516 6916 19572
rect 7644 24444 7700 24500
rect 7420 23436 7476 23492
rect 7420 23100 7476 23156
rect 7420 21868 7476 21924
rect 7532 21474 7588 21476
rect 7532 21422 7534 21474
rect 7534 21422 7586 21474
rect 7586 21422 7588 21474
rect 7532 21420 7588 21422
rect 9548 25282 9604 25284
rect 9548 25230 9550 25282
rect 9550 25230 9602 25282
rect 9602 25230 9604 25282
rect 9548 25228 9604 25230
rect 7868 23548 7924 23604
rect 7868 23042 7924 23044
rect 7868 22990 7870 23042
rect 7870 22990 7922 23042
rect 7922 22990 7924 23042
rect 7868 22988 7924 22990
rect 9548 24444 9604 24500
rect 9996 24220 10052 24276
rect 8652 24050 8708 24052
rect 8652 23998 8654 24050
rect 8654 23998 8706 24050
rect 8706 23998 8708 24050
rect 8652 23996 8708 23998
rect 8316 23826 8372 23828
rect 8316 23774 8318 23826
rect 8318 23774 8370 23826
rect 8370 23774 8372 23826
rect 8316 23772 8372 23774
rect 8092 22876 8148 22932
rect 8204 23100 8260 23156
rect 7644 20972 7700 21028
rect 8092 21532 8148 21588
rect 7756 20636 7812 20692
rect 7980 20690 8036 20692
rect 7980 20638 7982 20690
rect 7982 20638 8034 20690
rect 8034 20638 8036 20690
rect 7980 20636 8036 20638
rect 7644 20578 7700 20580
rect 7644 20526 7646 20578
rect 7646 20526 7698 20578
rect 7698 20526 7700 20578
rect 7644 20524 7700 20526
rect 8540 22876 8596 22932
rect 8540 22146 8596 22148
rect 8540 22094 8542 22146
rect 8542 22094 8594 22146
rect 8594 22094 8596 22146
rect 8540 22092 8596 22094
rect 7868 20076 7924 20132
rect 7084 19740 7140 19796
rect 7196 19906 7252 19908
rect 7196 19854 7198 19906
rect 7198 19854 7250 19906
rect 7250 19854 7252 19906
rect 7196 19852 7252 19854
rect 7084 19346 7140 19348
rect 7084 19294 7086 19346
rect 7086 19294 7138 19346
rect 7138 19294 7140 19346
rect 7084 19292 7140 19294
rect 6972 17164 7028 17220
rect 7196 17948 7252 18004
rect 7196 17666 7252 17668
rect 7196 17614 7198 17666
rect 7198 17614 7250 17666
rect 7250 17614 7252 17666
rect 7196 17612 7252 17614
rect 7644 19122 7700 19124
rect 7644 19070 7646 19122
rect 7646 19070 7698 19122
rect 7698 19070 7700 19122
rect 7644 19068 7700 19070
rect 7532 18284 7588 18340
rect 7532 17666 7588 17668
rect 7532 17614 7534 17666
rect 7534 17614 7586 17666
rect 7586 17614 7588 17666
rect 7532 17612 7588 17614
rect 7420 17442 7476 17444
rect 7420 17390 7422 17442
rect 7422 17390 7474 17442
rect 7474 17390 7476 17442
rect 7420 17388 7476 17390
rect 6860 16044 6916 16100
rect 6748 15932 6804 15988
rect 7308 16044 7364 16100
rect 7084 15874 7140 15876
rect 7084 15822 7086 15874
rect 7086 15822 7138 15874
rect 7138 15822 7140 15874
rect 7084 15820 7140 15822
rect 7308 15596 7364 15652
rect 7420 15484 7476 15540
rect 7756 16268 7812 16324
rect 8316 21196 8372 21252
rect 8092 19404 8148 19460
rect 8540 20578 8596 20580
rect 8540 20526 8542 20578
rect 8542 20526 8594 20578
rect 8594 20526 8596 20578
rect 8540 20524 8596 20526
rect 8540 20018 8596 20020
rect 8540 19966 8542 20018
rect 8542 19966 8594 20018
rect 8594 19966 8596 20018
rect 8540 19964 8596 19966
rect 8204 19292 8260 19348
rect 8316 19404 8372 19460
rect 8092 19122 8148 19124
rect 8092 19070 8094 19122
rect 8094 19070 8146 19122
rect 8146 19070 8148 19122
rect 8092 19068 8148 19070
rect 8092 18620 8148 18676
rect 7980 18172 8036 18228
rect 8316 18620 8372 18676
rect 8540 18508 8596 18564
rect 9100 24050 9156 24052
rect 9100 23998 9102 24050
rect 9102 23998 9154 24050
rect 9154 23998 9156 24050
rect 9100 23996 9156 23998
rect 8764 23436 8820 23492
rect 8764 22092 8820 22148
rect 9660 23548 9716 23604
rect 9100 21756 9156 21812
rect 9212 22204 9268 22260
rect 8988 20914 9044 20916
rect 8988 20862 8990 20914
rect 8990 20862 9042 20914
rect 9042 20862 9044 20914
rect 8988 20860 9044 20862
rect 9100 20524 9156 20580
rect 11116 24610 11172 24612
rect 11116 24558 11118 24610
rect 11118 24558 11170 24610
rect 11170 24558 11172 24610
rect 11116 24556 11172 24558
rect 11228 24332 11284 24388
rect 11564 24332 11620 24388
rect 11452 23884 11508 23940
rect 10892 23548 10948 23604
rect 10668 23212 10724 23268
rect 10220 23154 10276 23156
rect 10220 23102 10222 23154
rect 10222 23102 10274 23154
rect 10274 23102 10276 23154
rect 10220 23100 10276 23102
rect 9996 22316 10052 22372
rect 10668 22876 10724 22932
rect 10108 22258 10164 22260
rect 10108 22206 10110 22258
rect 10110 22206 10162 22258
rect 10162 22206 10164 22258
rect 10108 22204 10164 22206
rect 9548 21644 9604 21700
rect 9772 21868 9828 21924
rect 8876 19740 8932 19796
rect 9324 20524 9380 20580
rect 8764 19404 8820 19460
rect 9212 19964 9268 20020
rect 8428 17890 8484 17892
rect 8428 17838 8430 17890
rect 8430 17838 8482 17890
rect 8482 17838 8484 17890
rect 8428 17836 8484 17838
rect 8204 17612 8260 17668
rect 8540 17554 8596 17556
rect 8540 17502 8542 17554
rect 8542 17502 8594 17554
rect 8594 17502 8596 17554
rect 8540 17500 8596 17502
rect 8428 17164 8484 17220
rect 8540 17052 8596 17108
rect 8316 16940 8372 16996
rect 8204 16882 8260 16884
rect 8204 16830 8206 16882
rect 8206 16830 8258 16882
rect 8258 16830 8260 16882
rect 8204 16828 8260 16830
rect 8092 16604 8148 16660
rect 6412 14252 6468 14308
rect 7084 15148 7140 15204
rect 6636 14140 6692 14196
rect 5964 12962 6020 12964
rect 5964 12910 5966 12962
rect 5966 12910 6018 12962
rect 6018 12910 6020 12962
rect 5964 12908 6020 12910
rect 5852 11676 5908 11732
rect 5740 11394 5796 11396
rect 5740 11342 5742 11394
rect 5742 11342 5794 11394
rect 5794 11342 5796 11394
rect 5740 11340 5796 11342
rect 5628 10722 5684 10724
rect 5628 10670 5630 10722
rect 5630 10670 5682 10722
rect 5682 10670 5684 10722
rect 5628 10668 5684 10670
rect 5740 10556 5796 10612
rect 6412 13522 6468 13524
rect 6412 13470 6414 13522
rect 6414 13470 6466 13522
rect 6466 13470 6468 13522
rect 6412 13468 6468 13470
rect 6748 14028 6804 14084
rect 7532 15202 7588 15204
rect 7532 15150 7534 15202
rect 7534 15150 7586 15202
rect 7586 15150 7588 15202
rect 7532 15148 7588 15150
rect 7644 15036 7700 15092
rect 7756 15820 7812 15876
rect 7420 14364 7476 14420
rect 7196 14252 7252 14308
rect 6412 12572 6468 12628
rect 6860 13132 6916 13188
rect 6300 12066 6356 12068
rect 6300 12014 6302 12066
rect 6302 12014 6354 12066
rect 6354 12014 6356 12066
rect 6300 12012 6356 12014
rect 6188 11564 6244 11620
rect 6748 12684 6804 12740
rect 7308 13858 7364 13860
rect 7308 13806 7310 13858
rect 7310 13806 7362 13858
rect 7362 13806 7364 13858
rect 7308 13804 7364 13806
rect 7196 13020 7252 13076
rect 6972 12850 7028 12852
rect 6972 12798 6974 12850
rect 6974 12798 7026 12850
rect 7026 12798 7028 12850
rect 6972 12796 7028 12798
rect 6748 11788 6804 11844
rect 6076 10780 6132 10836
rect 6188 10610 6244 10612
rect 6188 10558 6190 10610
rect 6190 10558 6242 10610
rect 6242 10558 6244 10610
rect 6188 10556 6244 10558
rect 6636 11394 6692 11396
rect 6636 11342 6638 11394
rect 6638 11342 6690 11394
rect 6690 11342 6692 11394
rect 6636 11340 6692 11342
rect 6524 10780 6580 10836
rect 6188 10332 6244 10388
rect 5740 9548 5796 9604
rect 5852 9042 5908 9044
rect 5852 8990 5854 9042
rect 5854 8990 5906 9042
rect 5906 8990 5908 9042
rect 5852 8988 5908 8990
rect 5964 8540 6020 8596
rect 6636 11004 6692 11060
rect 7308 13580 7364 13636
rect 8988 18956 9044 19012
rect 9100 19292 9156 19348
rect 9436 19964 9492 20020
rect 9212 17388 9268 17444
rect 9100 17106 9156 17108
rect 9100 17054 9102 17106
rect 9102 17054 9154 17106
rect 9154 17054 9156 17106
rect 9100 17052 9156 17054
rect 8764 16940 8820 16996
rect 8652 16716 8708 16772
rect 8652 16380 8708 16436
rect 8204 15260 8260 15316
rect 7980 14700 8036 14756
rect 7868 14028 7924 14084
rect 8540 15148 8596 15204
rect 8092 14306 8148 14308
rect 8092 14254 8094 14306
rect 8094 14254 8146 14306
rect 8146 14254 8148 14306
rect 8092 14252 8148 14254
rect 8988 16268 9044 16324
rect 8764 15484 8820 15540
rect 8988 15260 9044 15316
rect 8764 14924 8820 14980
rect 8652 14252 8708 14308
rect 8876 13970 8932 13972
rect 8876 13918 8878 13970
rect 8878 13918 8930 13970
rect 8930 13918 8932 13970
rect 8876 13916 8932 13918
rect 8204 13858 8260 13860
rect 8204 13806 8206 13858
rect 8206 13806 8258 13858
rect 8258 13806 8260 13858
rect 8204 13804 8260 13806
rect 8764 13858 8820 13860
rect 8764 13806 8766 13858
rect 8766 13806 8818 13858
rect 8818 13806 8820 13858
rect 8764 13804 8820 13806
rect 7868 13746 7924 13748
rect 7868 13694 7870 13746
rect 7870 13694 7922 13746
rect 7922 13694 7924 13746
rect 7868 13692 7924 13694
rect 8204 13074 8260 13076
rect 8204 13022 8206 13074
rect 8206 13022 8258 13074
rect 8258 13022 8260 13074
rect 8204 13020 8260 13022
rect 7420 12738 7476 12740
rect 7420 12686 7422 12738
rect 7422 12686 7474 12738
rect 7474 12686 7476 12738
rect 7420 12684 7476 12686
rect 7532 12572 7588 12628
rect 8092 12684 8148 12740
rect 7196 12460 7252 12516
rect 7532 12348 7588 12404
rect 6972 11788 7028 11844
rect 7196 11676 7252 11732
rect 6860 10892 6916 10948
rect 6748 10498 6804 10500
rect 6748 10446 6750 10498
rect 6750 10446 6802 10498
rect 6802 10446 6804 10498
rect 6748 10444 6804 10446
rect 6412 9548 6468 9604
rect 6524 9436 6580 9492
rect 6524 9266 6580 9268
rect 6524 9214 6526 9266
rect 6526 9214 6578 9266
rect 6578 9214 6580 9266
rect 6524 9212 6580 9214
rect 6412 9154 6468 9156
rect 6412 9102 6414 9154
rect 6414 9102 6466 9154
rect 6466 9102 6468 9154
rect 6412 9100 6468 9102
rect 6300 9042 6356 9044
rect 6300 8990 6302 9042
rect 6302 8990 6354 9042
rect 6354 8990 6356 9042
rect 6300 8988 6356 8990
rect 7756 12236 7812 12292
rect 7532 11116 7588 11172
rect 7644 11788 7700 11844
rect 7308 10668 7364 10724
rect 7084 9996 7140 10052
rect 9100 13132 9156 13188
rect 8428 12962 8484 12964
rect 8428 12910 8430 12962
rect 8430 12910 8482 12962
rect 8482 12910 8484 12962
rect 8428 12908 8484 12910
rect 8876 12796 8932 12852
rect 8988 12572 9044 12628
rect 8316 11676 8372 11732
rect 7420 10556 7476 10612
rect 7196 9324 7252 9380
rect 7084 9266 7140 9268
rect 7084 9214 7086 9266
rect 7086 9214 7138 9266
rect 7138 9214 7140 9266
rect 7084 9212 7140 9214
rect 7532 10444 7588 10500
rect 7756 9996 7812 10052
rect 7644 9826 7700 9828
rect 7644 9774 7646 9826
rect 7646 9774 7698 9826
rect 7698 9774 7700 9826
rect 7644 9772 7700 9774
rect 7980 9772 8036 9828
rect 8092 9884 8148 9940
rect 7532 9154 7588 9156
rect 7532 9102 7534 9154
rect 7534 9102 7586 9154
rect 7586 9102 7588 9154
rect 7532 9100 7588 9102
rect 6860 8428 6916 8484
rect 6300 8258 6356 8260
rect 6300 8206 6302 8258
rect 6302 8206 6354 8258
rect 6354 8206 6356 8258
rect 6300 8204 6356 8206
rect 5628 8034 5684 8036
rect 5628 7982 5630 8034
rect 5630 7982 5682 8034
rect 5682 7982 5684 8034
rect 5628 7980 5684 7982
rect 4732 7474 4788 7476
rect 4732 7422 4734 7474
rect 4734 7422 4786 7474
rect 4786 7422 4788 7474
rect 4732 7420 4788 7422
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4620 6860 4676 6916
rect 4732 6690 4788 6692
rect 4732 6638 4734 6690
rect 4734 6638 4786 6690
rect 4786 6638 4788 6690
rect 4732 6636 4788 6638
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 5516 7474 5572 7476
rect 5516 7422 5518 7474
rect 5518 7422 5570 7474
rect 5570 7422 5572 7474
rect 5516 7420 5572 7422
rect 5068 6748 5124 6804
rect 5068 5964 5124 6020
rect 4956 5234 5012 5236
rect 4956 5182 4958 5234
rect 4958 5182 5010 5234
rect 5010 5182 5012 5234
rect 4956 5180 5012 5182
rect 4732 4732 4788 4788
rect 4844 4956 4900 5012
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4956 4060 5012 4116
rect 5180 5852 5236 5908
rect 5964 7362 6020 7364
rect 5964 7310 5966 7362
rect 5966 7310 6018 7362
rect 6018 7310 6020 7362
rect 5964 7308 6020 7310
rect 5628 6636 5684 6692
rect 6636 7980 6692 8036
rect 6524 7644 6580 7700
rect 5964 7084 6020 7140
rect 6076 6748 6132 6804
rect 5628 6466 5684 6468
rect 5628 6414 5630 6466
rect 5630 6414 5682 6466
rect 5682 6414 5684 6466
rect 5628 6412 5684 6414
rect 5516 6018 5572 6020
rect 5516 5966 5518 6018
rect 5518 5966 5570 6018
rect 5570 5966 5572 6018
rect 5516 5964 5572 5966
rect 5404 5404 5460 5460
rect 5852 5346 5908 5348
rect 5852 5294 5854 5346
rect 5854 5294 5906 5346
rect 5906 5294 5908 5346
rect 5852 5292 5908 5294
rect 5628 5180 5684 5236
rect 5852 5068 5908 5124
rect 6188 5964 6244 6020
rect 6412 7084 6468 7140
rect 6860 7644 6916 7700
rect 7084 8876 7140 8932
rect 7308 7698 7364 7700
rect 7308 7646 7310 7698
rect 7310 7646 7362 7698
rect 7362 7646 7364 7698
rect 7308 7644 7364 7646
rect 6636 7532 6692 7588
rect 6860 7474 6916 7476
rect 6860 7422 6862 7474
rect 6862 7422 6914 7474
rect 6914 7422 6916 7474
rect 6860 7420 6916 7422
rect 6748 7308 6804 7364
rect 6860 6636 6916 6692
rect 7308 7420 7364 7476
rect 7756 9324 7812 9380
rect 7868 9436 7924 9492
rect 7644 8034 7700 8036
rect 7644 7982 7646 8034
rect 7646 7982 7698 8034
rect 7698 7982 7700 8034
rect 7644 7980 7700 7982
rect 7644 7196 7700 7252
rect 7532 6524 7588 6580
rect 7308 6188 7364 6244
rect 6972 5740 7028 5796
rect 6860 5068 6916 5124
rect 6636 4844 6692 4900
rect 6188 4620 6244 4676
rect 6524 4450 6580 4452
rect 6524 4398 6526 4450
rect 6526 4398 6578 4450
rect 6578 4398 6580 4450
rect 6524 4396 6580 4398
rect 6188 3724 6244 3780
rect 7644 5068 7700 5124
rect 7420 4844 7476 4900
rect 6972 4562 7028 4564
rect 6972 4510 6974 4562
rect 6974 4510 7026 4562
rect 7026 4510 7028 4562
rect 6972 4508 7028 4510
rect 7644 4450 7700 4452
rect 7644 4398 7646 4450
rect 7646 4398 7698 4450
rect 7698 4398 7700 4450
rect 7644 4396 7700 4398
rect 6860 4284 6916 4340
rect 6748 3666 6804 3668
rect 6748 3614 6750 3666
rect 6750 3614 6802 3666
rect 6802 3614 6804 3666
rect 6748 3612 6804 3614
rect 3836 2604 3892 2660
rect 6412 3330 6468 3332
rect 6412 3278 6414 3330
rect 6414 3278 6466 3330
rect 6466 3278 6468 3330
rect 6412 3276 6468 3278
rect 7980 7586 8036 7588
rect 7980 7534 7982 7586
rect 7982 7534 8034 7586
rect 8034 7534 8036 7586
rect 7980 7532 8036 7534
rect 8428 10834 8484 10836
rect 8428 10782 8430 10834
rect 8430 10782 8482 10834
rect 8482 10782 8484 10834
rect 8428 10780 8484 10782
rect 8316 10332 8372 10388
rect 8540 10108 8596 10164
rect 8764 11900 8820 11956
rect 8204 9548 8260 9604
rect 8428 9436 8484 9492
rect 8204 8818 8260 8820
rect 8204 8766 8206 8818
rect 8206 8766 8258 8818
rect 8258 8766 8260 8818
rect 8204 8764 8260 8766
rect 8204 8428 8260 8484
rect 9100 12402 9156 12404
rect 9100 12350 9102 12402
rect 9102 12350 9154 12402
rect 9154 12350 9156 12402
rect 9100 12348 9156 12350
rect 9436 19740 9492 19796
rect 9436 18396 9492 18452
rect 9884 20412 9940 20468
rect 9660 19740 9716 19796
rect 9884 19180 9940 19236
rect 9884 18674 9940 18676
rect 9884 18622 9886 18674
rect 9886 18622 9938 18674
rect 9938 18622 9940 18674
rect 9884 18620 9940 18622
rect 9772 18562 9828 18564
rect 9772 18510 9774 18562
rect 9774 18510 9826 18562
rect 9826 18510 9828 18562
rect 9772 18508 9828 18510
rect 9660 17948 9716 18004
rect 9660 17388 9716 17444
rect 9436 16380 9492 16436
rect 9660 16604 9716 16660
rect 9324 16268 9380 16324
rect 9548 16156 9604 16212
rect 9324 15484 9380 15540
rect 9548 15484 9604 15540
rect 9324 14700 9380 14756
rect 9324 11788 9380 11844
rect 9324 11618 9380 11620
rect 9324 11566 9326 11618
rect 9326 11566 9378 11618
rect 9378 11566 9380 11618
rect 9324 11564 9380 11566
rect 9212 11452 9268 11508
rect 8876 11394 8932 11396
rect 8876 11342 8878 11394
rect 8878 11342 8930 11394
rect 8930 11342 8932 11394
rect 8876 11340 8932 11342
rect 9100 10780 9156 10836
rect 9324 11004 9380 11060
rect 9884 18226 9940 18228
rect 9884 18174 9886 18226
rect 9886 18174 9938 18226
rect 9938 18174 9940 18226
rect 9884 18172 9940 18174
rect 9772 14700 9828 14756
rect 10444 22146 10500 22148
rect 10444 22094 10446 22146
rect 10446 22094 10498 22146
rect 10498 22094 10500 22146
rect 10444 22092 10500 22094
rect 10668 21980 10724 22036
rect 10108 21810 10164 21812
rect 10108 21758 10110 21810
rect 10110 21758 10162 21810
rect 10162 21758 10164 21810
rect 10108 21756 10164 21758
rect 10556 21810 10612 21812
rect 10556 21758 10558 21810
rect 10558 21758 10610 21810
rect 10610 21758 10612 21810
rect 10556 21756 10612 21758
rect 10668 21644 10724 21700
rect 10220 20578 10276 20580
rect 10220 20526 10222 20578
rect 10222 20526 10274 20578
rect 10274 20526 10276 20578
rect 10220 20524 10276 20526
rect 10668 20188 10724 20244
rect 10444 20018 10500 20020
rect 10444 19966 10446 20018
rect 10446 19966 10498 20018
rect 10498 19966 10500 20018
rect 10444 19964 10500 19966
rect 10444 19234 10500 19236
rect 10444 19182 10446 19234
rect 10446 19182 10498 19234
rect 10498 19182 10500 19234
rect 10444 19180 10500 19182
rect 9884 17500 9940 17556
rect 10108 19068 10164 19124
rect 9660 14252 9716 14308
rect 9996 15484 10052 15540
rect 10668 19068 10724 19124
rect 11004 21868 11060 21924
rect 10892 20130 10948 20132
rect 10892 20078 10894 20130
rect 10894 20078 10946 20130
rect 10946 20078 10948 20130
rect 10892 20076 10948 20078
rect 10892 19852 10948 19908
rect 10332 17612 10388 17668
rect 10220 16994 10276 16996
rect 10220 16942 10222 16994
rect 10222 16942 10274 16994
rect 10274 16942 10276 16994
rect 10220 16940 10276 16942
rect 10556 16882 10612 16884
rect 10556 16830 10558 16882
rect 10558 16830 10610 16882
rect 10610 16830 10612 16882
rect 10556 16828 10612 16830
rect 9884 13916 9940 13972
rect 9996 14924 10052 14980
rect 10332 15708 10388 15764
rect 10556 15484 10612 15540
rect 10444 15260 10500 15316
rect 10332 15148 10388 15204
rect 10220 13970 10276 13972
rect 10220 13918 10222 13970
rect 10222 13918 10274 13970
rect 10274 13918 10276 13970
rect 10220 13916 10276 13918
rect 10108 13804 10164 13860
rect 9884 13356 9940 13412
rect 9772 11788 9828 11844
rect 9996 11788 10052 11844
rect 9884 11676 9940 11732
rect 9772 11452 9828 11508
rect 9772 11116 9828 11172
rect 8988 10108 9044 10164
rect 8540 8876 8596 8932
rect 8540 8428 8596 8484
rect 8876 8428 8932 8484
rect 8988 8764 9044 8820
rect 8316 8316 8372 8372
rect 8316 7980 8372 8036
rect 7980 7084 8036 7140
rect 8764 8034 8820 8036
rect 8764 7982 8766 8034
rect 8766 7982 8818 8034
rect 8818 7982 8820 8034
rect 8764 7980 8820 7982
rect 8428 7756 8484 7812
rect 8876 7644 8932 7700
rect 8652 7250 8708 7252
rect 8652 7198 8654 7250
rect 8654 7198 8706 7250
rect 8706 7198 8708 7250
rect 8652 7196 8708 7198
rect 8092 6188 8148 6244
rect 7868 3724 7924 3780
rect 7868 3442 7924 3444
rect 7868 3390 7870 3442
rect 7870 3390 7922 3442
rect 7922 3390 7924 3442
rect 7868 3388 7924 3390
rect 8876 6188 8932 6244
rect 8428 4956 8484 5012
rect 9100 7698 9156 7700
rect 9100 7646 9102 7698
rect 9102 7646 9154 7698
rect 9154 7646 9156 7698
rect 9100 7644 9156 7646
rect 9772 10610 9828 10612
rect 9772 10558 9774 10610
rect 9774 10558 9826 10610
rect 9826 10558 9828 10610
rect 9772 10556 9828 10558
rect 9772 9826 9828 9828
rect 9772 9774 9774 9826
rect 9774 9774 9826 9826
rect 9826 9774 9828 9826
rect 9772 9772 9828 9774
rect 9548 9714 9604 9716
rect 9548 9662 9550 9714
rect 9550 9662 9602 9714
rect 9602 9662 9604 9714
rect 9548 9660 9604 9662
rect 9996 11116 10052 11172
rect 10220 13356 10276 13412
rect 10220 12684 10276 12740
rect 10220 11788 10276 11844
rect 10220 11452 10276 11508
rect 9996 10780 10052 10836
rect 10892 18674 10948 18676
rect 10892 18622 10894 18674
rect 10894 18622 10946 18674
rect 10946 18622 10948 18674
rect 10892 18620 10948 18622
rect 11004 18562 11060 18564
rect 11004 18510 11006 18562
rect 11006 18510 11058 18562
rect 11058 18510 11060 18562
rect 11004 18508 11060 18510
rect 10892 18226 10948 18228
rect 10892 18174 10894 18226
rect 10894 18174 10946 18226
rect 10946 18174 10948 18226
rect 10892 18172 10948 18174
rect 11340 22482 11396 22484
rect 11340 22430 11342 22482
rect 11342 22430 11394 22482
rect 11394 22430 11396 22482
rect 11340 22428 11396 22430
rect 12236 24050 12292 24052
rect 12236 23998 12238 24050
rect 12238 23998 12290 24050
rect 12290 23998 12292 24050
rect 12236 23996 12292 23998
rect 14476 24332 14532 24388
rect 13468 23996 13524 24052
rect 14028 24108 14084 24164
rect 15036 24050 15092 24052
rect 15036 23998 15038 24050
rect 15038 23998 15090 24050
rect 15090 23998 15092 24050
rect 15036 23996 15092 23998
rect 13580 23938 13636 23940
rect 13580 23886 13582 23938
rect 13582 23886 13634 23938
rect 13634 23886 13636 23938
rect 13580 23884 13636 23886
rect 11564 20860 11620 20916
rect 11340 20242 11396 20244
rect 11340 20190 11342 20242
rect 11342 20190 11394 20242
rect 11394 20190 11396 20242
rect 11340 20188 11396 20190
rect 11228 18620 11284 18676
rect 11228 17554 11284 17556
rect 11228 17502 11230 17554
rect 11230 17502 11282 17554
rect 11282 17502 11284 17554
rect 11228 17500 11284 17502
rect 10892 16716 10948 16772
rect 10892 15260 10948 15316
rect 10780 14924 10836 14980
rect 10892 13916 10948 13972
rect 11228 16828 11284 16884
rect 11340 16604 11396 16660
rect 11676 23548 11732 23604
rect 11900 23548 11956 23604
rect 12684 23714 12740 23716
rect 12684 23662 12686 23714
rect 12686 23662 12738 23714
rect 12738 23662 12740 23714
rect 12684 23660 12740 23662
rect 11788 21756 11844 21812
rect 12012 21474 12068 21476
rect 12012 21422 12014 21474
rect 12014 21422 12066 21474
rect 12066 21422 12068 21474
rect 12012 21420 12068 21422
rect 11900 20914 11956 20916
rect 11900 20862 11902 20914
rect 11902 20862 11954 20914
rect 11954 20862 11956 20914
rect 11900 20860 11956 20862
rect 12124 20748 12180 20804
rect 12236 22764 12292 22820
rect 11676 19404 11732 19460
rect 12012 19906 12068 19908
rect 12012 19854 12014 19906
rect 12014 19854 12066 19906
rect 12066 19854 12068 19906
rect 12012 19852 12068 19854
rect 11788 18732 11844 18788
rect 12348 22146 12404 22148
rect 12348 22094 12350 22146
rect 12350 22094 12402 22146
rect 12402 22094 12404 22146
rect 12348 22092 12404 22094
rect 12348 21868 12404 21924
rect 13020 23154 13076 23156
rect 13020 23102 13022 23154
rect 13022 23102 13074 23154
rect 13074 23102 13076 23154
rect 13020 23100 13076 23102
rect 14028 23100 14084 23156
rect 12684 22988 12740 23044
rect 13804 23042 13860 23044
rect 13804 22990 13806 23042
rect 13806 22990 13858 23042
rect 13858 22990 13860 23042
rect 13804 22988 13860 22990
rect 13468 22876 13524 22932
rect 14028 22204 14084 22260
rect 12684 22092 12740 22148
rect 12908 21868 12964 21924
rect 13132 22092 13188 22148
rect 12908 20748 12964 20804
rect 12460 20578 12516 20580
rect 12460 20526 12462 20578
rect 12462 20526 12514 20578
rect 12514 20526 12516 20578
rect 12460 20524 12516 20526
rect 12908 20188 12964 20244
rect 12460 20130 12516 20132
rect 12460 20078 12462 20130
rect 12462 20078 12514 20130
rect 12514 20078 12516 20130
rect 12460 20076 12516 20078
rect 12348 19964 12404 20020
rect 12572 19404 12628 19460
rect 11900 18508 11956 18564
rect 12012 18956 12068 19012
rect 11452 18172 11508 18228
rect 12236 18508 12292 18564
rect 11676 17500 11732 17556
rect 11564 17164 11620 17220
rect 11900 16994 11956 16996
rect 11900 16942 11902 16994
rect 11902 16942 11954 16994
rect 11954 16942 11956 16994
rect 11900 16940 11956 16942
rect 11788 16882 11844 16884
rect 11788 16830 11790 16882
rect 11790 16830 11842 16882
rect 11842 16830 11844 16882
rect 11788 16828 11844 16830
rect 12124 17612 12180 17668
rect 12124 16716 12180 16772
rect 12236 16604 12292 16660
rect 11452 15986 11508 15988
rect 11452 15934 11454 15986
rect 11454 15934 11506 15986
rect 11506 15934 11508 15986
rect 11452 15932 11508 15934
rect 11116 15708 11172 15764
rect 11116 15314 11172 15316
rect 11116 15262 11118 15314
rect 11118 15262 11170 15314
rect 11170 15262 11172 15314
rect 11116 15260 11172 15262
rect 11564 15314 11620 15316
rect 11564 15262 11566 15314
rect 11566 15262 11618 15314
rect 11618 15262 11620 15314
rect 11564 15260 11620 15262
rect 11676 14700 11732 14756
rect 12348 18172 12404 18228
rect 12124 16156 12180 16212
rect 11900 15986 11956 15988
rect 11900 15934 11902 15986
rect 11902 15934 11954 15986
rect 11954 15934 11956 15986
rect 11900 15932 11956 15934
rect 12012 15874 12068 15876
rect 12012 15822 12014 15874
rect 12014 15822 12066 15874
rect 12066 15822 12068 15874
rect 12012 15820 12068 15822
rect 11900 15538 11956 15540
rect 11900 15486 11902 15538
rect 11902 15486 11954 15538
rect 11954 15486 11956 15538
rect 11900 15484 11956 15486
rect 11788 15036 11844 15092
rect 11228 14252 11284 14308
rect 12124 15372 12180 15428
rect 11116 14028 11172 14084
rect 11788 14252 11844 14308
rect 12012 14028 12068 14084
rect 11564 13468 11620 13524
rect 12460 17612 12516 17668
rect 12684 19010 12740 19012
rect 12684 18958 12686 19010
rect 12686 18958 12738 19010
rect 12738 18958 12740 19010
rect 12684 18956 12740 18958
rect 12684 18732 12740 18788
rect 12908 18284 12964 18340
rect 12796 18226 12852 18228
rect 12796 18174 12798 18226
rect 12798 18174 12850 18226
rect 12850 18174 12852 18226
rect 12796 18172 12852 18174
rect 13020 17948 13076 18004
rect 12684 17666 12740 17668
rect 12684 17614 12686 17666
rect 12686 17614 12738 17666
rect 12738 17614 12740 17666
rect 12684 17612 12740 17614
rect 12908 17500 12964 17556
rect 12684 17164 12740 17220
rect 12796 17388 12852 17444
rect 12796 16716 12852 16772
rect 12572 16604 12628 16660
rect 12684 16492 12740 16548
rect 12796 16322 12852 16324
rect 12796 16270 12798 16322
rect 12798 16270 12850 16322
rect 12850 16270 12852 16322
rect 12796 16268 12852 16270
rect 12684 15708 12740 15764
rect 12796 15986 12852 15988
rect 12796 15934 12798 15986
rect 12798 15934 12850 15986
rect 12850 15934 12852 15986
rect 12796 15932 12852 15934
rect 12572 15596 12628 15652
rect 12908 15708 12964 15764
rect 12684 15260 12740 15316
rect 12460 15202 12516 15204
rect 12460 15150 12462 15202
rect 12462 15150 12514 15202
rect 12514 15150 12516 15202
rect 12460 15148 12516 15150
rect 12572 14364 12628 14420
rect 12460 13916 12516 13972
rect 13020 15372 13076 15428
rect 12796 13858 12852 13860
rect 12796 13806 12798 13858
rect 12798 13806 12850 13858
rect 12850 13806 12852 13858
rect 12796 13804 12852 13806
rect 11004 12290 11060 12292
rect 11004 12238 11006 12290
rect 11006 12238 11058 12290
rect 11058 12238 11060 12290
rect 11004 12236 11060 12238
rect 10668 11564 10724 11620
rect 10220 10386 10276 10388
rect 10220 10334 10222 10386
rect 10222 10334 10274 10386
rect 10274 10334 10276 10386
rect 10220 10332 10276 10334
rect 11004 10780 11060 10836
rect 10780 10332 10836 10388
rect 10220 10108 10276 10164
rect 9996 9602 10052 9604
rect 9996 9550 9998 9602
rect 9998 9550 10050 9602
rect 10050 9550 10052 9602
rect 9996 9548 10052 9550
rect 11564 12236 11620 12292
rect 11228 11394 11284 11396
rect 11228 11342 11230 11394
rect 11230 11342 11282 11394
rect 11282 11342 11284 11394
rect 11228 11340 11284 11342
rect 11452 11340 11508 11396
rect 11228 10610 11284 10612
rect 11228 10558 11230 10610
rect 11230 10558 11282 10610
rect 11282 10558 11284 10610
rect 11228 10556 11284 10558
rect 11340 10386 11396 10388
rect 11340 10334 11342 10386
rect 11342 10334 11394 10386
rect 11394 10334 11396 10386
rect 11340 10332 11396 10334
rect 10780 9714 10836 9716
rect 10780 9662 10782 9714
rect 10782 9662 10834 9714
rect 10834 9662 10836 9714
rect 10780 9660 10836 9662
rect 9324 7196 9380 7252
rect 9548 8764 9604 8820
rect 8988 4956 9044 5012
rect 8988 4620 9044 4676
rect 9324 6972 9380 7028
rect 10108 8988 10164 9044
rect 9996 8258 10052 8260
rect 9996 8206 9998 8258
rect 9998 8206 10050 8258
rect 10050 8206 10052 8258
rect 9996 8204 10052 8206
rect 9884 7644 9940 7700
rect 9772 6860 9828 6916
rect 9996 7196 10052 7252
rect 9996 6412 10052 6468
rect 9884 6076 9940 6132
rect 10444 8876 10500 8932
rect 10780 8764 10836 8820
rect 10892 9602 10948 9604
rect 10892 9550 10894 9602
rect 10894 9550 10946 9602
rect 10946 9550 10948 9602
rect 10892 9548 10948 9550
rect 10892 8652 10948 8708
rect 10444 8540 10500 8596
rect 10332 8428 10388 8484
rect 10556 7474 10612 7476
rect 10556 7422 10558 7474
rect 10558 7422 10610 7474
rect 10610 7422 10612 7474
rect 10556 7420 10612 7422
rect 10780 7698 10836 7700
rect 10780 7646 10782 7698
rect 10782 7646 10834 7698
rect 10834 7646 10836 7698
rect 10780 7644 10836 7646
rect 11228 8652 11284 8708
rect 11004 7196 11060 7252
rect 11228 8204 11284 8260
rect 10556 7084 10612 7140
rect 11228 6748 11284 6804
rect 9212 5628 9268 5684
rect 9884 4732 9940 4788
rect 9772 4620 9828 4676
rect 9100 4172 9156 4228
rect 9212 4396 9268 4452
rect 8876 3724 8932 3780
rect 7196 3164 7252 3220
rect 7084 2716 7140 2772
rect 10220 5740 10276 5796
rect 11004 5292 11060 5348
rect 9996 4060 10052 4116
rect 10108 5068 10164 5124
rect 10556 4396 10612 4452
rect 11228 4396 11284 4452
rect 12460 13468 12516 13524
rect 12684 13468 12740 13524
rect 11676 12012 11732 12068
rect 12236 11788 12292 11844
rect 12572 12012 12628 12068
rect 12572 11228 12628 11284
rect 11676 11170 11732 11172
rect 11676 11118 11678 11170
rect 11678 11118 11730 11170
rect 11730 11118 11732 11170
rect 11676 11116 11732 11118
rect 12460 11170 12516 11172
rect 12460 11118 12462 11170
rect 12462 11118 12514 11170
rect 12514 11118 12516 11170
rect 12460 11116 12516 11118
rect 11564 10444 11620 10500
rect 11900 10498 11956 10500
rect 11900 10446 11902 10498
rect 11902 10446 11954 10498
rect 11954 10446 11956 10498
rect 11900 10444 11956 10446
rect 12124 9772 12180 9828
rect 11564 7980 11620 8036
rect 12012 7532 12068 7588
rect 12236 9154 12292 9156
rect 12236 9102 12238 9154
rect 12238 9102 12290 9154
rect 12290 9102 12292 9154
rect 12236 9100 12292 9102
rect 12796 9884 12852 9940
rect 12684 9714 12740 9716
rect 12684 9662 12686 9714
rect 12686 9662 12738 9714
rect 12738 9662 12740 9714
rect 12684 9660 12740 9662
rect 12796 9324 12852 9380
rect 13020 9602 13076 9604
rect 13020 9550 13022 9602
rect 13022 9550 13074 9602
rect 13074 9550 13076 9602
rect 13020 9548 13076 9550
rect 12908 8540 12964 8596
rect 14140 22146 14196 22148
rect 14140 22094 14142 22146
rect 14142 22094 14194 22146
rect 14194 22094 14196 22146
rect 14140 22092 14196 22094
rect 14140 21868 14196 21924
rect 15148 22204 15204 22260
rect 14700 21532 14756 21588
rect 15372 22146 15428 22148
rect 15372 22094 15374 22146
rect 15374 22094 15426 22146
rect 15426 22094 15428 22146
rect 15372 22092 15428 22094
rect 15484 21868 15540 21924
rect 14924 21644 14980 21700
rect 14476 21196 14532 21252
rect 14476 20972 14532 21028
rect 13356 20130 13412 20132
rect 13356 20078 13358 20130
rect 13358 20078 13410 20130
rect 13410 20078 13412 20130
rect 13356 20076 13412 20078
rect 13244 18508 13300 18564
rect 14924 20972 14980 21028
rect 15372 21420 15428 21476
rect 14028 19906 14084 19908
rect 14028 19854 14030 19906
rect 14030 19854 14082 19906
rect 14082 19854 14084 19906
rect 14028 19852 14084 19854
rect 13580 19404 13636 19460
rect 14252 19404 14308 19460
rect 14140 19010 14196 19012
rect 14140 18958 14142 19010
rect 14142 18958 14194 19010
rect 14194 18958 14196 19010
rect 14140 18956 14196 18958
rect 14252 18620 14308 18676
rect 13468 18396 13524 18452
rect 14028 18508 14084 18564
rect 13356 17724 13412 17780
rect 13804 17442 13860 17444
rect 13804 17390 13806 17442
rect 13806 17390 13858 17442
rect 13858 17390 13860 17442
rect 13804 17388 13860 17390
rect 13580 17106 13636 17108
rect 13580 17054 13582 17106
rect 13582 17054 13634 17106
rect 13634 17054 13636 17106
rect 13580 17052 13636 17054
rect 13692 16828 13748 16884
rect 13804 16268 13860 16324
rect 14140 17724 14196 17780
rect 14140 17276 14196 17332
rect 14028 17164 14084 17220
rect 15036 20130 15092 20132
rect 15036 20078 15038 20130
rect 15038 20078 15090 20130
rect 15090 20078 15092 20130
rect 15036 20076 15092 20078
rect 14588 18956 14644 19012
rect 14700 18508 14756 18564
rect 14476 17612 14532 17668
rect 14588 18396 14644 18452
rect 14812 18284 14868 18340
rect 14924 18956 14980 19012
rect 14476 17388 14532 17444
rect 15036 18508 15092 18564
rect 15148 17948 15204 18004
rect 14252 17052 14308 17108
rect 14476 17164 14532 17220
rect 14028 16940 14084 16996
rect 13468 15932 13524 15988
rect 13692 16098 13748 16100
rect 13692 16046 13694 16098
rect 13694 16046 13746 16098
rect 13746 16046 13748 16098
rect 13692 16044 13748 16046
rect 13356 15484 13412 15540
rect 13804 15932 13860 15988
rect 13692 15260 13748 15316
rect 13468 15036 13524 15092
rect 13468 14588 13524 14644
rect 13916 15874 13972 15876
rect 13916 15822 13918 15874
rect 13918 15822 13970 15874
rect 13970 15822 13972 15874
rect 13916 15820 13972 15822
rect 14252 16604 14308 16660
rect 14140 16492 14196 16548
rect 14588 17052 14644 17108
rect 14700 16828 14756 16884
rect 14476 16492 14532 16548
rect 14812 16604 14868 16660
rect 14924 16268 14980 16324
rect 14140 14588 14196 14644
rect 13244 14140 13300 14196
rect 14028 14530 14084 14532
rect 14028 14478 14030 14530
rect 14030 14478 14082 14530
rect 14082 14478 14084 14530
rect 14028 14476 14084 14478
rect 13356 13692 13412 13748
rect 14588 15986 14644 15988
rect 14588 15934 14590 15986
rect 14590 15934 14642 15986
rect 14642 15934 14644 15986
rect 14588 15932 14644 15934
rect 14812 16044 14868 16100
rect 14812 15708 14868 15764
rect 14924 15932 14980 15988
rect 14588 15596 14644 15652
rect 14588 15314 14644 15316
rect 14588 15262 14590 15314
rect 14590 15262 14642 15314
rect 14642 15262 14644 15314
rect 14588 15260 14644 15262
rect 14700 15484 14756 15540
rect 14476 14924 14532 14980
rect 15484 19516 15540 19572
rect 15372 17836 15428 17892
rect 15708 18620 15764 18676
rect 15372 17666 15428 17668
rect 15372 17614 15374 17666
rect 15374 17614 15426 17666
rect 15426 17614 15428 17666
rect 15372 17612 15428 17614
rect 15372 16940 15428 16996
rect 15260 16716 15316 16772
rect 15596 18338 15652 18340
rect 15596 18286 15598 18338
rect 15598 18286 15650 18338
rect 15650 18286 15652 18338
rect 15596 18284 15652 18286
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 20972 25228 21028 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19516 24220 19572 24276
rect 19404 23996 19460 24052
rect 17612 23772 17668 23828
rect 16828 23154 16884 23156
rect 16828 23102 16830 23154
rect 16830 23102 16882 23154
rect 16882 23102 16884 23154
rect 16828 23100 16884 23102
rect 16940 22988 16996 23044
rect 16492 22764 16548 22820
rect 16828 22764 16884 22820
rect 16044 22316 16100 22372
rect 16492 22258 16548 22260
rect 16492 22206 16494 22258
rect 16494 22206 16546 22258
rect 16546 22206 16548 22258
rect 16492 22204 16548 22206
rect 16156 22146 16212 22148
rect 16156 22094 16158 22146
rect 16158 22094 16210 22146
rect 16210 22094 16212 22146
rect 16156 22092 16212 22094
rect 16156 21868 16212 21924
rect 17388 22482 17444 22484
rect 17388 22430 17390 22482
rect 17390 22430 17442 22482
rect 17442 22430 17444 22482
rect 17388 22428 17444 22430
rect 16940 22146 16996 22148
rect 16940 22094 16942 22146
rect 16942 22094 16994 22146
rect 16994 22094 16996 22146
rect 16940 22092 16996 22094
rect 17836 22540 17892 22596
rect 17612 21810 17668 21812
rect 17612 21758 17614 21810
rect 17614 21758 17666 21810
rect 17666 21758 17668 21810
rect 17612 21756 17668 21758
rect 16044 21698 16100 21700
rect 16044 21646 16046 21698
rect 16046 21646 16098 21698
rect 16098 21646 16100 21698
rect 16044 21644 16100 21646
rect 16492 21698 16548 21700
rect 16492 21646 16494 21698
rect 16494 21646 16546 21698
rect 16546 21646 16548 21698
rect 18060 22204 18116 22260
rect 16492 21644 16548 21646
rect 15932 20076 15988 20132
rect 16156 21532 16212 21588
rect 16268 20578 16324 20580
rect 16268 20526 16270 20578
rect 16270 20526 16322 20578
rect 16322 20526 16324 20578
rect 16268 20524 16324 20526
rect 16156 20300 16212 20356
rect 15820 18172 15876 18228
rect 16044 18956 16100 19012
rect 16604 20188 16660 20244
rect 16940 20524 16996 20580
rect 16716 19906 16772 19908
rect 16716 19854 16718 19906
rect 16718 19854 16770 19906
rect 16770 19854 16772 19906
rect 16716 19852 16772 19854
rect 17948 20578 18004 20580
rect 17948 20526 17950 20578
rect 17950 20526 18002 20578
rect 18002 20526 18004 20578
rect 17948 20524 18004 20526
rect 17388 20300 17444 20356
rect 16940 19740 16996 19796
rect 16380 18956 16436 19012
rect 15596 16828 15652 16884
rect 15708 17948 15764 18004
rect 16156 17948 16212 18004
rect 15932 17164 15988 17220
rect 16044 16940 16100 16996
rect 16156 17052 16212 17108
rect 15148 15708 15204 15764
rect 15372 15986 15428 15988
rect 15372 15934 15374 15986
rect 15374 15934 15426 15986
rect 15426 15934 15428 15986
rect 15372 15932 15428 15934
rect 15036 14700 15092 14756
rect 14812 14642 14868 14644
rect 14812 14590 14814 14642
rect 14814 14590 14866 14642
rect 14866 14590 14868 14642
rect 14812 14588 14868 14590
rect 15036 14530 15092 14532
rect 15036 14478 15038 14530
rect 15038 14478 15090 14530
rect 15090 14478 15092 14530
rect 15036 14476 15092 14478
rect 14588 14364 14644 14420
rect 15260 15314 15316 15316
rect 15260 15262 15262 15314
rect 15262 15262 15314 15314
rect 15314 15262 15316 15314
rect 15260 15260 15316 15262
rect 15148 13916 15204 13972
rect 15260 14140 15316 14196
rect 14476 13522 14532 13524
rect 14476 13470 14478 13522
rect 14478 13470 14530 13522
rect 14530 13470 14532 13522
rect 14476 13468 14532 13470
rect 14812 13468 14868 13524
rect 14924 13580 14980 13636
rect 14364 13186 14420 13188
rect 14364 13134 14366 13186
rect 14366 13134 14418 13186
rect 14418 13134 14420 13186
rect 14364 13132 14420 13134
rect 15036 13244 15092 13300
rect 14588 13020 14644 13076
rect 13692 12850 13748 12852
rect 13692 12798 13694 12850
rect 13694 12798 13746 12850
rect 13746 12798 13748 12850
rect 13692 12796 13748 12798
rect 13356 9996 13412 10052
rect 13692 9826 13748 9828
rect 13692 9774 13694 9826
rect 13694 9774 13746 9826
rect 13746 9774 13748 9826
rect 13692 9772 13748 9774
rect 14028 11116 14084 11172
rect 14812 12962 14868 12964
rect 14812 12910 14814 12962
rect 14814 12910 14866 12962
rect 14866 12910 14868 12962
rect 14812 12908 14868 12910
rect 14588 12348 14644 12404
rect 14588 12066 14644 12068
rect 14588 12014 14590 12066
rect 14590 12014 14642 12066
rect 14642 12014 14644 12066
rect 14588 12012 14644 12014
rect 14924 11564 14980 11620
rect 14700 11282 14756 11284
rect 14700 11230 14702 11282
rect 14702 11230 14754 11282
rect 14754 11230 14756 11282
rect 14700 11228 14756 11230
rect 14812 10780 14868 10836
rect 14252 10108 14308 10164
rect 14924 10444 14980 10500
rect 14140 9996 14196 10052
rect 13916 9826 13972 9828
rect 13916 9774 13918 9826
rect 13918 9774 13970 9826
rect 13970 9774 13972 9826
rect 13916 9772 13972 9774
rect 13468 9266 13524 9268
rect 13468 9214 13470 9266
rect 13470 9214 13522 9266
rect 13522 9214 13524 9266
rect 13468 9212 13524 9214
rect 13132 8204 13188 8260
rect 12684 7644 12740 7700
rect 12348 6748 12404 6804
rect 11564 6018 11620 6020
rect 11564 5966 11566 6018
rect 11566 5966 11618 6018
rect 11618 5966 11620 6018
rect 11564 5964 11620 5966
rect 11452 5740 11508 5796
rect 10332 4172 10388 4228
rect 11228 4060 11284 4116
rect 10668 3836 10724 3892
rect 10556 3778 10612 3780
rect 10556 3726 10558 3778
rect 10558 3726 10610 3778
rect 10610 3726 10612 3778
rect 10556 3724 10612 3726
rect 11900 5404 11956 5460
rect 13580 8930 13636 8932
rect 13580 8878 13582 8930
rect 13582 8878 13634 8930
rect 13634 8878 13636 8930
rect 13580 8876 13636 8878
rect 14252 9884 14308 9940
rect 13692 8316 13748 8372
rect 13804 8540 13860 8596
rect 13692 8146 13748 8148
rect 13692 8094 13694 8146
rect 13694 8094 13746 8146
rect 13746 8094 13748 8146
rect 13692 8092 13748 8094
rect 14140 8204 14196 8260
rect 14140 7980 14196 8036
rect 13804 6636 13860 6692
rect 12460 6578 12516 6580
rect 12460 6526 12462 6578
rect 12462 6526 12514 6578
rect 12514 6526 12516 6578
rect 12460 6524 12516 6526
rect 12012 4508 12068 4564
rect 11452 3836 11508 3892
rect 11676 3500 11732 3556
rect 12572 5122 12628 5124
rect 12572 5070 12574 5122
rect 12574 5070 12626 5122
rect 12626 5070 12628 5122
rect 12572 5068 12628 5070
rect 12348 5010 12404 5012
rect 12348 4958 12350 5010
rect 12350 4958 12402 5010
rect 12402 4958 12404 5010
rect 12348 4956 12404 4958
rect 12796 6466 12852 6468
rect 12796 6414 12798 6466
rect 12798 6414 12850 6466
rect 12850 6414 12852 6466
rect 12796 6412 12852 6414
rect 14140 6578 14196 6580
rect 14140 6526 14142 6578
rect 14142 6526 14194 6578
rect 14194 6526 14196 6578
rect 14140 6524 14196 6526
rect 13916 6300 13972 6356
rect 14476 7756 14532 7812
rect 14588 9436 14644 9492
rect 14924 9884 14980 9940
rect 15036 9772 15092 9828
rect 14700 9324 14756 9380
rect 14588 6524 14644 6580
rect 14364 6188 14420 6244
rect 13468 5794 13524 5796
rect 13468 5742 13470 5794
rect 13470 5742 13522 5794
rect 13522 5742 13524 5794
rect 13468 5740 13524 5742
rect 12684 4284 12740 4340
rect 13916 4396 13972 4452
rect 16268 16882 16324 16884
rect 16268 16830 16270 16882
rect 16270 16830 16322 16882
rect 16322 16830 16324 16882
rect 16268 16828 16324 16830
rect 16492 17836 16548 17892
rect 16492 17106 16548 17108
rect 16492 17054 16494 17106
rect 16494 17054 16546 17106
rect 16546 17054 16548 17106
rect 16492 17052 16548 17054
rect 17612 19852 17668 19908
rect 17388 19010 17444 19012
rect 17388 18958 17390 19010
rect 17390 18958 17442 19010
rect 17442 18958 17444 19010
rect 17388 18956 17444 18958
rect 16940 18844 16996 18900
rect 17052 18508 17108 18564
rect 16828 17836 16884 17892
rect 16604 16882 16660 16884
rect 16604 16830 16606 16882
rect 16606 16830 16658 16882
rect 16658 16830 16660 16882
rect 16604 16828 16660 16830
rect 16940 16940 16996 16996
rect 15820 16044 15876 16100
rect 15708 15986 15764 15988
rect 15708 15934 15710 15986
rect 15710 15934 15762 15986
rect 15762 15934 15764 15986
rect 15708 15932 15764 15934
rect 15708 15708 15764 15764
rect 15820 15148 15876 15204
rect 16380 15708 16436 15764
rect 16492 15484 16548 15540
rect 16156 15148 16212 15204
rect 15932 14588 15988 14644
rect 16268 14530 16324 14532
rect 16268 14478 16270 14530
rect 16270 14478 16322 14530
rect 16322 14478 16324 14530
rect 16268 14476 16324 14478
rect 15596 13746 15652 13748
rect 15596 13694 15598 13746
rect 15598 13694 15650 13746
rect 15650 13694 15652 13746
rect 15596 13692 15652 13694
rect 15372 13468 15428 13524
rect 15372 11564 15428 11620
rect 15372 10780 15428 10836
rect 15820 13858 15876 13860
rect 15820 13806 15822 13858
rect 15822 13806 15874 13858
rect 15874 13806 15876 13858
rect 15820 13804 15876 13806
rect 15820 13468 15876 13524
rect 16828 15484 16884 15540
rect 17836 19292 17892 19348
rect 17612 18508 17668 18564
rect 17388 18172 17444 18228
rect 18284 22146 18340 22148
rect 18284 22094 18286 22146
rect 18286 22094 18338 22146
rect 18338 22094 18340 22146
rect 18284 22092 18340 22094
rect 18284 21868 18340 21924
rect 18172 21474 18228 21476
rect 18172 21422 18174 21474
rect 18174 21422 18226 21474
rect 18226 21422 18228 21474
rect 18172 21420 18228 21422
rect 18508 21474 18564 21476
rect 18508 21422 18510 21474
rect 18510 21422 18562 21474
rect 18562 21422 18564 21474
rect 18508 21420 18564 21422
rect 18732 20578 18788 20580
rect 18732 20526 18734 20578
rect 18734 20526 18786 20578
rect 18786 20526 18788 20578
rect 18732 20524 18788 20526
rect 18060 19346 18116 19348
rect 18060 19294 18062 19346
rect 18062 19294 18114 19346
rect 18114 19294 18116 19346
rect 18060 19292 18116 19294
rect 18172 20076 18228 20132
rect 17388 16940 17444 16996
rect 18060 18620 18116 18676
rect 18508 19122 18564 19124
rect 18508 19070 18510 19122
rect 18510 19070 18562 19122
rect 18562 19070 18564 19122
rect 18508 19068 18564 19070
rect 18620 19516 18676 19572
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 18956 19122 19012 19124
rect 18956 19070 18958 19122
rect 18958 19070 19010 19122
rect 19010 19070 19012 19122
rect 18956 19068 19012 19070
rect 17724 16994 17780 16996
rect 17724 16942 17726 16994
rect 17726 16942 17778 16994
rect 17778 16942 17780 16994
rect 17724 16940 17780 16942
rect 18508 17164 18564 17220
rect 18508 16994 18564 16996
rect 18508 16942 18510 16994
rect 18510 16942 18562 16994
rect 18562 16942 18564 16994
rect 18508 16940 18564 16942
rect 17164 15986 17220 15988
rect 17164 15934 17166 15986
rect 17166 15934 17218 15986
rect 17218 15934 17220 15986
rect 17164 15932 17220 15934
rect 17164 15596 17220 15652
rect 16716 14140 16772 14196
rect 16604 13916 16660 13972
rect 15596 12572 15652 12628
rect 15820 12460 15876 12516
rect 15708 11228 15764 11284
rect 16268 12572 16324 12628
rect 16268 12236 16324 12292
rect 16268 11340 16324 11396
rect 16156 11282 16212 11284
rect 16156 11230 16158 11282
rect 16158 11230 16210 11282
rect 16210 11230 16212 11282
rect 16156 11228 16212 11230
rect 15820 10892 15876 10948
rect 16156 10780 16212 10836
rect 15596 9996 15652 10052
rect 16044 9938 16100 9940
rect 16044 9886 16046 9938
rect 16046 9886 16098 9938
rect 16098 9886 16100 9938
rect 16044 9884 16100 9886
rect 15260 9772 15316 9828
rect 16716 13746 16772 13748
rect 16716 13694 16718 13746
rect 16718 13694 16770 13746
rect 16770 13694 16772 13746
rect 16716 13692 16772 13694
rect 16828 13132 16884 13188
rect 17276 15372 17332 15428
rect 17276 14306 17332 14308
rect 17276 14254 17278 14306
rect 17278 14254 17330 14306
rect 17330 14254 17332 14306
rect 17276 14252 17332 14254
rect 17052 14140 17108 14196
rect 17388 13132 17444 13188
rect 17948 16098 18004 16100
rect 17948 16046 17950 16098
rect 17950 16046 18002 16098
rect 18002 16046 18004 16098
rect 17948 16044 18004 16046
rect 17836 15538 17892 15540
rect 17836 15486 17838 15538
rect 17838 15486 17890 15538
rect 17890 15486 17892 15538
rect 17836 15484 17892 15486
rect 17948 15314 18004 15316
rect 17948 15262 17950 15314
rect 17950 15262 18002 15314
rect 18002 15262 18004 15314
rect 17948 15260 18004 15262
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20300 21756 20356 21812
rect 19628 20690 19684 20692
rect 19628 20638 19630 20690
rect 19630 20638 19682 20690
rect 19682 20638 19684 20690
rect 19628 20636 19684 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19852 20188 19908 20244
rect 19292 19906 19348 19908
rect 19292 19854 19294 19906
rect 19294 19854 19346 19906
rect 19346 19854 19348 19906
rect 19292 19852 19348 19854
rect 19404 19346 19460 19348
rect 19404 19294 19406 19346
rect 19406 19294 19458 19346
rect 19458 19294 19460 19346
rect 19404 19292 19460 19294
rect 19180 18508 19236 18564
rect 20076 19906 20132 19908
rect 20076 19854 20078 19906
rect 20078 19854 20130 19906
rect 20130 19854 20132 19906
rect 20076 19852 20132 19854
rect 19852 19010 19908 19012
rect 19852 18958 19854 19010
rect 19854 18958 19906 19010
rect 19906 18958 19908 19010
rect 19852 18956 19908 18958
rect 19068 18396 19124 18452
rect 18732 17106 18788 17108
rect 18732 17054 18734 17106
rect 18734 17054 18786 17106
rect 18786 17054 18788 17106
rect 18732 17052 18788 17054
rect 18844 16322 18900 16324
rect 18844 16270 18846 16322
rect 18846 16270 18898 16322
rect 18898 16270 18900 16322
rect 18844 16268 18900 16270
rect 18732 15986 18788 15988
rect 18732 15934 18734 15986
rect 18734 15934 18786 15986
rect 18786 15934 18788 15986
rect 18732 15932 18788 15934
rect 18284 15874 18340 15876
rect 18284 15822 18286 15874
rect 18286 15822 18338 15874
rect 18338 15822 18340 15874
rect 18284 15820 18340 15822
rect 18844 15820 18900 15876
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20524 20860 20580 20916
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 42700 23884 42756 23940
rect 21308 23100 21364 23156
rect 20300 19346 20356 19348
rect 20300 19294 20302 19346
rect 20302 19294 20354 19346
rect 20354 19294 20356 19346
rect 20300 19292 20356 19294
rect 19068 17500 19124 17556
rect 19180 18338 19236 18340
rect 19180 18286 19182 18338
rect 19182 18286 19234 18338
rect 19234 18286 19236 18338
rect 19180 18284 19236 18286
rect 19068 16994 19124 16996
rect 19068 16942 19070 16994
rect 19070 16942 19122 16994
rect 19122 16942 19124 16994
rect 19068 16940 19124 16942
rect 19068 15932 19124 15988
rect 18396 15372 18452 15428
rect 17836 14252 17892 14308
rect 16940 12572 16996 12628
rect 16492 11116 16548 11172
rect 16380 10556 16436 10612
rect 16940 12348 16996 12404
rect 16604 10444 16660 10500
rect 16268 10332 16324 10388
rect 15148 9436 15204 9492
rect 16492 9772 16548 9828
rect 15148 8764 15204 8820
rect 15484 9042 15540 9044
rect 15484 8990 15486 9042
rect 15486 8990 15538 9042
rect 15538 8990 15540 9042
rect 15484 8988 15540 8990
rect 14812 8092 14868 8148
rect 15260 7756 15316 7812
rect 15820 9042 15876 9044
rect 15820 8990 15822 9042
rect 15822 8990 15874 9042
rect 15874 8990 15876 9042
rect 15820 8988 15876 8990
rect 16492 9042 16548 9044
rect 16492 8990 16494 9042
rect 16494 8990 16546 9042
rect 16546 8990 16548 9042
rect 16492 8988 16548 8990
rect 15484 8540 15540 8596
rect 15820 8428 15876 8484
rect 15372 7644 15428 7700
rect 15596 8204 15652 8260
rect 16044 7868 16100 7924
rect 16380 7644 16436 7700
rect 16716 11900 16772 11956
rect 16828 11452 16884 11508
rect 16828 10108 16884 10164
rect 16828 9714 16884 9716
rect 16828 9662 16830 9714
rect 16830 9662 16882 9714
rect 16882 9662 16884 9714
rect 16828 9660 16884 9662
rect 17052 10722 17108 10724
rect 17052 10670 17054 10722
rect 17054 10670 17106 10722
rect 17106 10670 17108 10722
rect 17052 10668 17108 10670
rect 17500 11452 17556 11508
rect 17388 11394 17444 11396
rect 17388 11342 17390 11394
rect 17390 11342 17442 11394
rect 17442 11342 17444 11394
rect 17388 11340 17444 11342
rect 17500 11282 17556 11284
rect 17500 11230 17502 11282
rect 17502 11230 17554 11282
rect 17554 11230 17556 11282
rect 17500 11228 17556 11230
rect 17276 11116 17332 11172
rect 17612 11170 17668 11172
rect 17612 11118 17614 11170
rect 17614 11118 17666 11170
rect 17666 11118 17668 11170
rect 17612 11116 17668 11118
rect 18172 14306 18228 14308
rect 18172 14254 18174 14306
rect 18174 14254 18226 14306
rect 18226 14254 18228 14306
rect 18172 14252 18228 14254
rect 18060 14140 18116 14196
rect 18172 13580 18228 13636
rect 18060 13522 18116 13524
rect 18060 13470 18062 13522
rect 18062 13470 18114 13522
rect 18114 13470 18116 13522
rect 18060 13468 18116 13470
rect 17948 13132 18004 13188
rect 18172 12124 18228 12180
rect 18060 11564 18116 11620
rect 17836 11116 17892 11172
rect 17052 10108 17108 10164
rect 17948 10108 18004 10164
rect 17948 9884 18004 9940
rect 18060 10332 18116 10388
rect 17724 9826 17780 9828
rect 17724 9774 17726 9826
rect 17726 9774 17778 9826
rect 17778 9774 17780 9826
rect 17724 9772 17780 9774
rect 17836 9714 17892 9716
rect 17836 9662 17838 9714
rect 17838 9662 17890 9714
rect 17890 9662 17892 9714
rect 17836 9660 17892 9662
rect 17836 9266 17892 9268
rect 17836 9214 17838 9266
rect 17838 9214 17890 9266
rect 17890 9214 17892 9266
rect 17836 9212 17892 9214
rect 17612 9042 17668 9044
rect 17612 8990 17614 9042
rect 17614 8990 17666 9042
rect 17666 8990 17668 9042
rect 17612 8988 17668 8990
rect 16940 8146 16996 8148
rect 16940 8094 16942 8146
rect 16942 8094 16994 8146
rect 16994 8094 16996 8146
rect 16940 8092 16996 8094
rect 16828 7868 16884 7924
rect 15596 6914 15652 6916
rect 15596 6862 15598 6914
rect 15598 6862 15650 6914
rect 15650 6862 15652 6914
rect 15596 6860 15652 6862
rect 17164 7756 17220 7812
rect 16716 6748 16772 6804
rect 15260 6524 15316 6580
rect 14252 5404 14308 5460
rect 14364 4844 14420 4900
rect 14140 4620 14196 4676
rect 14812 5234 14868 5236
rect 14812 5182 14814 5234
rect 14814 5182 14866 5234
rect 14866 5182 14868 5234
rect 14812 5180 14868 5182
rect 12796 3666 12852 3668
rect 12796 3614 12798 3666
rect 12798 3614 12850 3666
rect 12850 3614 12852 3666
rect 12796 3612 12852 3614
rect 15372 6300 15428 6356
rect 15708 6188 15764 6244
rect 15820 6018 15876 6020
rect 15820 5966 15822 6018
rect 15822 5966 15874 6018
rect 15874 5966 15876 6018
rect 15820 5964 15876 5966
rect 16044 5180 16100 5236
rect 15148 4732 15204 4788
rect 14700 4338 14756 4340
rect 14700 4286 14702 4338
rect 14702 4286 14754 4338
rect 14754 4286 14756 4338
rect 14700 4284 14756 4286
rect 14028 3612 14084 3668
rect 14588 3666 14644 3668
rect 14588 3614 14590 3666
rect 14590 3614 14642 3666
rect 14642 3614 14644 3666
rect 14588 3612 14644 3614
rect 15484 3666 15540 3668
rect 15484 3614 15486 3666
rect 15486 3614 15538 3666
rect 15538 3614 15540 3666
rect 15484 3612 15540 3614
rect 10220 3052 10276 3108
rect 10556 3276 10612 3332
rect 13244 3500 13300 3556
rect 14700 3388 14756 3444
rect 13916 2940 13972 2996
rect 17052 6914 17108 6916
rect 17052 6862 17054 6914
rect 17054 6862 17106 6914
rect 17106 6862 17108 6914
rect 17052 6860 17108 6862
rect 16940 6466 16996 6468
rect 16940 6414 16942 6466
rect 16942 6414 16994 6466
rect 16994 6414 16996 6466
rect 16940 6412 16996 6414
rect 16828 6188 16884 6244
rect 16940 6130 16996 6132
rect 16940 6078 16942 6130
rect 16942 6078 16994 6130
rect 16994 6078 16996 6130
rect 16940 6076 16996 6078
rect 16828 6018 16884 6020
rect 16828 5966 16830 6018
rect 16830 5966 16882 6018
rect 16882 5966 16884 6018
rect 16828 5964 16884 5966
rect 16828 5628 16884 5684
rect 16716 5404 16772 5460
rect 17052 5292 17108 5348
rect 16716 4732 16772 4788
rect 16828 4396 16884 4452
rect 16492 3612 16548 3668
rect 17724 7698 17780 7700
rect 17724 7646 17726 7698
rect 17726 7646 17778 7698
rect 17778 7646 17780 7698
rect 17724 7644 17780 7646
rect 17500 7084 17556 7140
rect 17276 6300 17332 6356
rect 17388 6636 17444 6692
rect 17388 5852 17444 5908
rect 17948 7698 18004 7700
rect 17948 7646 17950 7698
rect 17950 7646 18002 7698
rect 18002 7646 18004 7698
rect 17948 7644 18004 7646
rect 18732 15314 18788 15316
rect 18732 15262 18734 15314
rect 18734 15262 18786 15314
rect 18786 15262 18788 15314
rect 18732 15260 18788 15262
rect 18508 14140 18564 14196
rect 18620 14924 18676 14980
rect 18956 15372 19012 15428
rect 18732 13916 18788 13972
rect 18844 13858 18900 13860
rect 18844 13806 18846 13858
rect 18846 13806 18898 13858
rect 18898 13806 18900 13858
rect 18844 13804 18900 13806
rect 18620 13692 18676 13748
rect 19292 17836 19348 17892
rect 20188 18338 20244 18340
rect 20188 18286 20190 18338
rect 20190 18286 20242 18338
rect 20242 18286 20244 18338
rect 20188 18284 20244 18286
rect 20300 17836 20356 17892
rect 19404 17442 19460 17444
rect 19404 17390 19406 17442
rect 19406 17390 19458 17442
rect 19458 17390 19460 17442
rect 19404 17388 19460 17390
rect 19964 17442 20020 17444
rect 19964 17390 19966 17442
rect 19966 17390 20018 17442
rect 20018 17390 20020 17442
rect 19964 17388 20020 17390
rect 19292 17276 19348 17332
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19180 15484 19236 15540
rect 19180 15148 19236 15204
rect 19516 16156 19572 16212
rect 19404 15986 19460 15988
rect 19404 15934 19406 15986
rect 19406 15934 19458 15986
rect 19458 15934 19460 15986
rect 19404 15932 19460 15934
rect 19516 15874 19572 15876
rect 19516 15822 19518 15874
rect 19518 15822 19570 15874
rect 19570 15822 19572 15874
rect 19516 15820 19572 15822
rect 20076 15932 20132 15988
rect 19740 15874 19796 15876
rect 19740 15822 19742 15874
rect 19742 15822 19794 15874
rect 19794 15822 19796 15874
rect 19740 15820 19796 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19628 15484 19684 15540
rect 19516 15148 19572 15204
rect 19404 14754 19460 14756
rect 19404 14702 19406 14754
rect 19406 14702 19458 14754
rect 19458 14702 19460 14754
rect 19404 14700 19460 14702
rect 20636 17388 20692 17444
rect 20860 17836 20916 17892
rect 20860 17164 20916 17220
rect 20636 16156 20692 16212
rect 20412 16098 20468 16100
rect 20412 16046 20414 16098
rect 20414 16046 20466 16098
rect 20466 16046 20468 16098
rect 20412 16044 20468 16046
rect 20860 16156 20916 16212
rect 20636 15596 20692 15652
rect 20748 15820 20804 15876
rect 20188 14700 20244 14756
rect 19516 14530 19572 14532
rect 19516 14478 19518 14530
rect 19518 14478 19570 14530
rect 19570 14478 19572 14530
rect 19516 14476 19572 14478
rect 20860 15538 20916 15540
rect 20860 15486 20862 15538
rect 20862 15486 20914 15538
rect 20914 15486 20916 15538
rect 20860 15484 20916 15486
rect 20412 15260 20468 15316
rect 20524 15036 20580 15092
rect 20076 14530 20132 14532
rect 20076 14478 20078 14530
rect 20078 14478 20130 14530
rect 20130 14478 20132 14530
rect 20076 14476 20132 14478
rect 20412 14476 20468 14532
rect 19292 14364 19348 14420
rect 19068 14028 19124 14084
rect 19404 14306 19460 14308
rect 19404 14254 19406 14306
rect 19406 14254 19458 14306
rect 19458 14254 19460 14306
rect 19404 14252 19460 14254
rect 19180 13692 19236 13748
rect 19068 13580 19124 13636
rect 18620 11564 18676 11620
rect 19836 14138 19892 14140
rect 19516 14028 19572 14084
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20636 14476 20692 14532
rect 20748 15260 20804 15316
rect 20300 14306 20356 14308
rect 20300 14254 20302 14306
rect 20302 14254 20354 14306
rect 20354 14254 20356 14306
rect 20300 14252 20356 14254
rect 20636 14306 20692 14308
rect 20636 14254 20638 14306
rect 20638 14254 20690 14306
rect 20690 14254 20692 14306
rect 20636 14252 20692 14254
rect 20412 14028 20468 14084
rect 20524 13804 20580 13860
rect 19628 13468 19684 13524
rect 19292 13356 19348 13412
rect 19852 13356 19908 13412
rect 19516 13244 19572 13300
rect 19068 12460 19124 12516
rect 18732 11170 18788 11172
rect 18732 11118 18734 11170
rect 18734 11118 18786 11170
rect 18786 11118 18788 11170
rect 18732 11116 18788 11118
rect 18620 11004 18676 11060
rect 18508 10780 18564 10836
rect 18508 10610 18564 10612
rect 18508 10558 18510 10610
rect 18510 10558 18562 10610
rect 18562 10558 18564 10610
rect 18508 10556 18564 10558
rect 18620 9884 18676 9940
rect 18956 9884 19012 9940
rect 18844 9548 18900 9604
rect 18396 8764 18452 8820
rect 19404 11394 19460 11396
rect 19404 11342 19406 11394
rect 19406 11342 19458 11394
rect 19458 11342 19460 11394
rect 19404 11340 19460 11342
rect 19292 10108 19348 10164
rect 19180 9772 19236 9828
rect 20076 12962 20132 12964
rect 20076 12910 20078 12962
rect 20078 12910 20130 12962
rect 20130 12910 20132 12962
rect 20076 12908 20132 12910
rect 19740 12850 19796 12852
rect 19740 12798 19742 12850
rect 19742 12798 19794 12850
rect 19794 12798 19796 12850
rect 19740 12796 19796 12798
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19628 12178 19684 12180
rect 19628 12126 19630 12178
rect 19630 12126 19682 12178
rect 19682 12126 19684 12178
rect 19628 12124 19684 12126
rect 20524 12236 20580 12292
rect 20412 11788 20468 11844
rect 21084 18338 21140 18340
rect 21084 18286 21086 18338
rect 21086 18286 21138 18338
rect 21138 18286 21140 18338
rect 21084 18284 21140 18286
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 42588 22540 42644 22596
rect 42252 22428 42308 22484
rect 25340 22316 25396 22372
rect 22316 22092 22372 22148
rect 21420 19740 21476 19796
rect 21532 17612 21588 17668
rect 21532 17276 21588 17332
rect 22540 20524 22596 20580
rect 22428 19628 22484 19684
rect 21868 18060 21924 18116
rect 21644 16828 21700 16884
rect 21756 17388 21812 17444
rect 21420 16268 21476 16324
rect 21644 16156 21700 16212
rect 21308 15820 21364 15876
rect 21532 15596 21588 15652
rect 21084 15260 21140 15316
rect 20860 13244 20916 13300
rect 21084 13244 21140 13300
rect 21868 16268 21924 16324
rect 21868 15314 21924 15316
rect 21868 15262 21870 15314
rect 21870 15262 21922 15314
rect 21922 15262 21924 15314
rect 21868 15260 21924 15262
rect 21756 14924 21812 14980
rect 21196 12908 21252 12964
rect 21420 13916 21476 13972
rect 23548 19292 23604 19348
rect 22876 18450 22932 18452
rect 22876 18398 22878 18450
rect 22878 18398 22930 18450
rect 22930 18398 22932 18450
rect 22876 18396 22932 18398
rect 22092 17442 22148 17444
rect 22092 17390 22094 17442
rect 22094 17390 22146 17442
rect 22146 17390 22148 17442
rect 22092 17388 22148 17390
rect 22652 18284 22708 18340
rect 23548 17778 23604 17780
rect 23548 17726 23550 17778
rect 23550 17726 23602 17778
rect 23602 17726 23604 17778
rect 23548 17724 23604 17726
rect 23100 17442 23156 17444
rect 23100 17390 23102 17442
rect 23102 17390 23154 17442
rect 23154 17390 23156 17442
rect 23100 17388 23156 17390
rect 22652 17106 22708 17108
rect 22652 17054 22654 17106
rect 22654 17054 22706 17106
rect 22706 17054 22708 17106
rect 22652 17052 22708 17054
rect 23548 17164 23604 17220
rect 22092 15484 22148 15540
rect 22204 15372 22260 15428
rect 22652 16716 22708 16772
rect 22764 16210 22820 16212
rect 22764 16158 22766 16210
rect 22766 16158 22818 16210
rect 22818 16158 22820 16210
rect 22764 16156 22820 16158
rect 22540 15314 22596 15316
rect 22540 15262 22542 15314
rect 22542 15262 22594 15314
rect 22594 15262 22596 15314
rect 22540 15260 22596 15262
rect 21980 14588 22036 14644
rect 21980 14418 22036 14420
rect 21980 14366 21982 14418
rect 21982 14366 22034 14418
rect 22034 14366 22036 14418
rect 21980 14364 22036 14366
rect 21756 14028 21812 14084
rect 21980 14028 22036 14084
rect 20860 12236 20916 12292
rect 19852 11170 19908 11172
rect 19852 11118 19854 11170
rect 19854 11118 19906 11170
rect 19906 11118 19908 11170
rect 19852 11116 19908 11118
rect 19628 11004 19684 11060
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19628 9884 19684 9940
rect 19516 9714 19572 9716
rect 19516 9662 19518 9714
rect 19518 9662 19570 9714
rect 19570 9662 19572 9714
rect 19516 9660 19572 9662
rect 19852 9714 19908 9716
rect 19852 9662 19854 9714
rect 19854 9662 19906 9714
rect 19906 9662 19908 9714
rect 19852 9660 19908 9662
rect 19740 9548 19796 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19404 8818 19460 8820
rect 19404 8766 19406 8818
rect 19406 8766 19458 8818
rect 19458 8766 19460 8818
rect 19404 8764 19460 8766
rect 19068 8540 19124 8596
rect 19292 8316 19348 8372
rect 18284 8092 18340 8148
rect 18284 7644 18340 7700
rect 18396 6412 18452 6468
rect 18396 5964 18452 6020
rect 18508 6524 18564 6580
rect 17724 5906 17780 5908
rect 17724 5854 17726 5906
rect 17726 5854 17778 5906
rect 17778 5854 17780 5906
rect 17724 5852 17780 5854
rect 18620 6300 18676 6356
rect 17500 4956 17556 5012
rect 18060 5068 18116 5124
rect 17164 3500 17220 3556
rect 17612 4620 17668 4676
rect 18284 4508 18340 4564
rect 18172 4338 18228 4340
rect 18172 4286 18174 4338
rect 18174 4286 18226 4338
rect 18226 4286 18228 4338
rect 18172 4284 18228 4286
rect 17724 3778 17780 3780
rect 17724 3726 17726 3778
rect 17726 3726 17778 3778
rect 17778 3726 17780 3778
rect 17724 3724 17780 3726
rect 17612 3554 17668 3556
rect 17612 3502 17614 3554
rect 17614 3502 17666 3554
rect 17666 3502 17668 3554
rect 17612 3500 17668 3502
rect 18508 5516 18564 5572
rect 18844 6690 18900 6692
rect 18844 6638 18846 6690
rect 18846 6638 18898 6690
rect 18898 6638 18900 6690
rect 18844 6636 18900 6638
rect 19292 7308 19348 7364
rect 19852 8988 19908 9044
rect 19852 8316 19908 8372
rect 20524 11116 20580 11172
rect 20524 10498 20580 10500
rect 20524 10446 20526 10498
rect 20526 10446 20578 10498
rect 20578 10446 20580 10498
rect 20524 10444 20580 10446
rect 20300 9548 20356 9604
rect 20412 9660 20468 9716
rect 20524 9602 20580 9604
rect 20524 9550 20526 9602
rect 20526 9550 20578 9602
rect 20578 9550 20580 9602
rect 20524 9548 20580 9550
rect 20636 9266 20692 9268
rect 20636 9214 20638 9266
rect 20638 9214 20690 9266
rect 20690 9214 20692 9266
rect 20636 9212 20692 9214
rect 20860 9996 20916 10052
rect 20860 9826 20916 9828
rect 20860 9774 20862 9826
rect 20862 9774 20914 9826
rect 20914 9774 20916 9826
rect 20860 9772 20916 9774
rect 20860 8876 20916 8932
rect 19740 7980 19796 8036
rect 19852 8092 19908 8148
rect 20300 7980 20356 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19628 7474 19684 7476
rect 19628 7422 19630 7474
rect 19630 7422 19682 7474
rect 19682 7422 19684 7474
rect 19628 7420 19684 7422
rect 19180 6860 19236 6916
rect 19292 6578 19348 6580
rect 19292 6526 19294 6578
rect 19294 6526 19346 6578
rect 19346 6526 19348 6578
rect 19292 6524 19348 6526
rect 19516 7362 19572 7364
rect 19516 7310 19518 7362
rect 19518 7310 19570 7362
rect 19570 7310 19572 7362
rect 19516 7308 19572 7310
rect 19404 6300 19460 6356
rect 19852 7420 19908 7476
rect 19068 6188 19124 6244
rect 19852 6972 19908 7028
rect 20188 7308 20244 7364
rect 20972 8428 21028 8484
rect 22204 14306 22260 14308
rect 22204 14254 22206 14306
rect 22206 14254 22258 14306
rect 22258 14254 22260 14306
rect 22204 14252 22260 14254
rect 22092 13916 22148 13972
rect 22764 15426 22820 15428
rect 22764 15374 22766 15426
rect 22766 15374 22818 15426
rect 22818 15374 22820 15426
rect 22764 15372 22820 15374
rect 22652 13804 22708 13860
rect 22764 14924 22820 14980
rect 22652 13634 22708 13636
rect 22652 13582 22654 13634
rect 22654 13582 22706 13634
rect 22706 13582 22708 13634
rect 22652 13580 22708 13582
rect 22988 14700 23044 14756
rect 22204 13468 22260 13524
rect 21420 11116 21476 11172
rect 21532 11340 21588 11396
rect 21084 9100 21140 9156
rect 21196 11004 21252 11060
rect 21420 9884 21476 9940
rect 21532 9772 21588 9828
rect 21644 12236 21700 12292
rect 21756 11900 21812 11956
rect 21980 12572 22036 12628
rect 21868 11788 21924 11844
rect 21420 9212 21476 9268
rect 21420 9042 21476 9044
rect 21420 8990 21422 9042
rect 21422 8990 21474 9042
rect 21474 8990 21476 9042
rect 21420 8988 21476 8990
rect 21420 8204 21476 8260
rect 20748 7644 20804 7700
rect 20524 7308 20580 7364
rect 20860 7474 20916 7476
rect 20860 7422 20862 7474
rect 20862 7422 20914 7474
rect 20914 7422 20916 7474
rect 20860 7420 20916 7422
rect 20636 6466 20692 6468
rect 20636 6414 20638 6466
rect 20638 6414 20690 6466
rect 20690 6414 20692 6466
rect 20636 6412 20692 6414
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20636 6076 20692 6132
rect 18508 3500 18564 3556
rect 15932 2940 15988 2996
rect 18732 3948 18788 4004
rect 19292 3948 19348 4004
rect 19516 3500 19572 3556
rect 20300 5628 20356 5684
rect 20300 5346 20356 5348
rect 20300 5294 20302 5346
rect 20302 5294 20354 5346
rect 20354 5294 20356 5346
rect 20300 5292 20356 5294
rect 19740 5068 19796 5124
rect 20524 5122 20580 5124
rect 20524 5070 20526 5122
rect 20526 5070 20578 5122
rect 20578 5070 20580 5122
rect 20524 5068 20580 5070
rect 20188 4956 20244 5012
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21868 11004 21924 11060
rect 21868 9996 21924 10052
rect 22764 13468 22820 13524
rect 22652 13356 22708 13412
rect 22540 13132 22596 13188
rect 22876 13244 22932 13300
rect 22316 12738 22372 12740
rect 22316 12686 22318 12738
rect 22318 12686 22370 12738
rect 22370 12686 22372 12738
rect 22316 12684 22372 12686
rect 22540 12460 22596 12516
rect 22316 12236 22372 12292
rect 22092 10668 22148 10724
rect 22204 11394 22260 11396
rect 22204 11342 22206 11394
rect 22206 11342 22258 11394
rect 22258 11342 22260 11394
rect 22204 11340 22260 11342
rect 22652 11788 22708 11844
rect 22764 12908 22820 12964
rect 22204 10556 22260 10612
rect 21980 9884 22036 9940
rect 21644 7980 21700 8036
rect 21532 7362 21588 7364
rect 21532 7310 21534 7362
rect 21534 7310 21586 7362
rect 21586 7310 21588 7362
rect 21532 7308 21588 7310
rect 21980 9602 22036 9604
rect 21980 9550 21982 9602
rect 21982 9550 22034 9602
rect 22034 9550 22036 9602
rect 21980 9548 22036 9550
rect 21980 8540 22036 8596
rect 21868 8146 21924 8148
rect 21868 8094 21870 8146
rect 21870 8094 21922 8146
rect 21922 8094 21924 8146
rect 21868 8092 21924 8094
rect 21756 6748 21812 6804
rect 22204 8428 22260 8484
rect 22092 7420 22148 7476
rect 21868 6636 21924 6692
rect 21644 6300 21700 6356
rect 21756 5964 21812 6020
rect 21868 5852 21924 5908
rect 21644 5404 21700 5460
rect 22764 11170 22820 11172
rect 22764 11118 22766 11170
rect 22766 11118 22818 11170
rect 22818 11118 22820 11170
rect 22764 11116 22820 11118
rect 22764 10332 22820 10388
rect 22652 9996 22708 10052
rect 23212 16210 23268 16212
rect 23212 16158 23214 16210
rect 23214 16158 23266 16210
rect 23266 16158 23268 16210
rect 23212 16156 23268 16158
rect 23212 15820 23268 15876
rect 23884 15372 23940 15428
rect 23212 15314 23268 15316
rect 23212 15262 23214 15314
rect 23214 15262 23266 15314
rect 23266 15262 23268 15314
rect 23212 15260 23268 15262
rect 23772 14924 23828 14980
rect 23996 14812 24052 14868
rect 23772 14700 23828 14756
rect 23324 13916 23380 13972
rect 23884 13804 23940 13860
rect 23100 12908 23156 12964
rect 23324 13468 23380 13524
rect 23548 13244 23604 13300
rect 23100 12684 23156 12740
rect 23772 12460 23828 12516
rect 23212 12402 23268 12404
rect 23212 12350 23214 12402
rect 23214 12350 23266 12402
rect 23266 12350 23268 12402
rect 23212 12348 23268 12350
rect 23492 12348 23548 12404
rect 22988 12124 23044 12180
rect 23436 12178 23492 12180
rect 23436 12126 23438 12178
rect 23438 12126 23490 12178
rect 23490 12126 23492 12178
rect 23436 12124 23492 12126
rect 23100 12012 23156 12068
rect 22988 9772 23044 9828
rect 23100 10444 23156 10500
rect 22764 8540 22820 8596
rect 22428 8316 22484 8372
rect 22428 7644 22484 7700
rect 23100 6860 23156 6916
rect 23324 12012 23380 12068
rect 23548 11676 23604 11732
rect 23660 12290 23716 12292
rect 23660 12238 23662 12290
rect 23662 12238 23714 12290
rect 23714 12238 23716 12290
rect 23660 12236 23716 12238
rect 23660 11564 23716 11620
rect 23996 12460 24052 12516
rect 24332 17106 24388 17108
rect 24332 17054 24334 17106
rect 24334 17054 24386 17106
rect 24386 17054 24388 17106
rect 24332 17052 24388 17054
rect 24780 16994 24836 16996
rect 24780 16942 24782 16994
rect 24782 16942 24834 16994
rect 24834 16942 24836 16994
rect 24780 16940 24836 16942
rect 24556 15484 24612 15540
rect 24444 15426 24500 15428
rect 24444 15374 24446 15426
rect 24446 15374 24498 15426
rect 24498 15374 24500 15426
rect 24444 15372 24500 15374
rect 25228 15874 25284 15876
rect 25228 15822 25230 15874
rect 25230 15822 25282 15874
rect 25282 15822 25284 15874
rect 25228 15820 25284 15822
rect 24892 15484 24948 15540
rect 24668 15372 24724 15428
rect 25228 15260 25284 15316
rect 24556 13970 24612 13972
rect 24556 13918 24558 13970
rect 24558 13918 24610 13970
rect 24610 13918 24612 13970
rect 24556 13916 24612 13918
rect 24444 13858 24500 13860
rect 24444 13806 24446 13858
rect 24446 13806 24498 13858
rect 24498 13806 24500 13858
rect 24444 13804 24500 13806
rect 24556 13522 24612 13524
rect 24556 13470 24558 13522
rect 24558 13470 24610 13522
rect 24610 13470 24612 13522
rect 24556 13468 24612 13470
rect 24332 13356 24388 13412
rect 24668 13356 24724 13412
rect 24220 13020 24276 13076
rect 24444 13074 24500 13076
rect 24444 13022 24446 13074
rect 24446 13022 24498 13074
rect 24498 13022 24500 13074
rect 24444 13020 24500 13022
rect 24108 12124 24164 12180
rect 24556 12684 24612 12740
rect 23884 11564 23940 11620
rect 23996 11394 24052 11396
rect 23996 11342 23998 11394
rect 23998 11342 24050 11394
rect 24050 11342 24052 11394
rect 23996 11340 24052 11342
rect 23548 9772 23604 9828
rect 23436 9212 23492 9268
rect 22428 6018 22484 6020
rect 22428 5966 22430 6018
rect 22430 5966 22482 6018
rect 22482 5966 22484 6018
rect 22428 5964 22484 5966
rect 22988 5852 23044 5908
rect 22204 5068 22260 5124
rect 22540 5068 22596 5124
rect 21644 4450 21700 4452
rect 21644 4398 21646 4450
rect 21646 4398 21698 4450
rect 21698 4398 21700 4450
rect 21644 4396 21700 4398
rect 21420 4060 21476 4116
rect 21532 3948 21588 4004
rect 22428 5010 22484 5012
rect 22428 4958 22430 5010
rect 22430 4958 22482 5010
rect 22482 4958 22484 5010
rect 22428 4956 22484 4958
rect 22092 4898 22148 4900
rect 22092 4846 22094 4898
rect 22094 4846 22146 4898
rect 22146 4846 22148 4898
rect 22092 4844 22148 4846
rect 22204 4396 22260 4452
rect 22316 4620 22372 4676
rect 21868 3836 21924 3892
rect 23212 5068 23268 5124
rect 23100 4732 23156 4788
rect 22988 4508 23044 4564
rect 23212 4508 23268 4564
rect 22316 3724 22372 3780
rect 17724 3164 17780 3220
rect 16828 2828 16884 2884
rect 17276 2828 17332 2884
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21308 3388 21364 3444
rect 22540 3442 22596 3444
rect 22540 3390 22542 3442
rect 22542 3390 22594 3442
rect 22594 3390 22596 3442
rect 22540 3388 22596 3390
rect 24444 11900 24500 11956
rect 24556 11676 24612 11732
rect 23884 10780 23940 10836
rect 23660 8988 23716 9044
rect 23772 9996 23828 10052
rect 23660 7362 23716 7364
rect 23660 7310 23662 7362
rect 23662 7310 23714 7362
rect 23714 7310 23716 7362
rect 23660 7308 23716 7310
rect 24556 10332 24612 10388
rect 24556 8764 24612 8820
rect 23884 8092 23940 8148
rect 24220 8540 24276 8596
rect 24444 7698 24500 7700
rect 24444 7646 24446 7698
rect 24446 7646 24498 7698
rect 24498 7646 24500 7698
rect 24444 7644 24500 7646
rect 24556 6972 24612 7028
rect 24220 6636 24276 6692
rect 24332 6860 24388 6916
rect 24220 6300 24276 6356
rect 24220 5906 24276 5908
rect 24220 5854 24222 5906
rect 24222 5854 24274 5906
rect 24274 5854 24276 5906
rect 24220 5852 24276 5854
rect 23548 3836 23604 3892
rect 23324 3388 23380 3444
rect 23996 5122 24052 5124
rect 23996 5070 23998 5122
rect 23998 5070 24050 5122
rect 24050 5070 24052 5122
rect 23996 5068 24052 5070
rect 24444 6130 24500 6132
rect 24444 6078 24446 6130
rect 24446 6078 24498 6130
rect 24498 6078 24500 6130
rect 24444 6076 24500 6078
rect 25004 12348 25060 12404
rect 24892 11788 24948 11844
rect 25116 11564 25172 11620
rect 25004 11340 25060 11396
rect 24892 11282 24948 11284
rect 24892 11230 24894 11282
rect 24894 11230 24946 11282
rect 24946 11230 24948 11282
rect 24892 11228 24948 11230
rect 25004 10220 25060 10276
rect 24892 9996 24948 10052
rect 39116 22370 39172 22372
rect 39116 22318 39118 22370
rect 39118 22318 39170 22370
rect 39170 22318 39172 22370
rect 39116 22316 39172 22318
rect 40572 22316 40628 22372
rect 40012 21980 40068 22036
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 26460 16882 26516 16884
rect 26460 16830 26462 16882
rect 26462 16830 26514 16882
rect 26514 16830 26516 16882
rect 26460 16828 26516 16830
rect 25676 15426 25732 15428
rect 25676 15374 25678 15426
rect 25678 15374 25730 15426
rect 25730 15374 25732 15426
rect 25676 15372 25732 15374
rect 25788 15202 25844 15204
rect 25788 15150 25790 15202
rect 25790 15150 25842 15202
rect 25842 15150 25844 15202
rect 25788 15148 25844 15150
rect 25452 14924 25508 14980
rect 25340 14812 25396 14868
rect 26124 15372 26180 15428
rect 26684 15260 26740 15316
rect 26012 15036 26068 15092
rect 25564 13804 25620 13860
rect 26012 14364 26068 14420
rect 26012 13746 26068 13748
rect 26012 13694 26014 13746
rect 26014 13694 26066 13746
rect 26066 13694 26068 13746
rect 26012 13692 26068 13694
rect 25564 13356 25620 13412
rect 25564 13186 25620 13188
rect 25564 13134 25566 13186
rect 25566 13134 25618 13186
rect 25618 13134 25620 13186
rect 25564 13132 25620 13134
rect 25676 12572 25732 12628
rect 25788 12402 25844 12404
rect 25788 12350 25790 12402
rect 25790 12350 25842 12402
rect 25842 12350 25844 12402
rect 25788 12348 25844 12350
rect 25340 11452 25396 11508
rect 25676 11676 25732 11732
rect 25788 11564 25844 11620
rect 26012 11394 26068 11396
rect 26012 11342 26014 11394
rect 26014 11342 26066 11394
rect 26066 11342 26068 11394
rect 26012 11340 26068 11342
rect 25900 11116 25956 11172
rect 25676 10108 25732 10164
rect 25788 10332 25844 10388
rect 25228 8876 25284 8932
rect 24892 8764 24948 8820
rect 24780 6412 24836 6468
rect 24892 8428 24948 8484
rect 25564 7868 25620 7924
rect 26348 13916 26404 13972
rect 26684 14306 26740 14308
rect 26684 14254 26686 14306
rect 26686 14254 26738 14306
rect 26738 14254 26740 14306
rect 26684 14252 26740 14254
rect 26572 13804 26628 13860
rect 26348 13468 26404 13524
rect 26460 12962 26516 12964
rect 26460 12910 26462 12962
rect 26462 12910 26514 12962
rect 26514 12910 26516 12962
rect 26460 12908 26516 12910
rect 26348 12460 26404 12516
rect 26684 13468 26740 13524
rect 26908 15148 26964 15204
rect 27132 15820 27188 15876
rect 27244 15260 27300 15316
rect 26796 13580 26852 13636
rect 26124 11116 26180 11172
rect 27132 14252 27188 14308
rect 27468 16770 27524 16772
rect 27468 16718 27470 16770
rect 27470 16718 27522 16770
rect 27522 16718 27524 16770
rect 27468 16716 27524 16718
rect 29484 16716 29540 16772
rect 27468 16492 27524 16548
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 29932 16210 29988 16212
rect 29932 16158 29934 16210
rect 29934 16158 29986 16210
rect 29986 16158 29988 16210
rect 29932 16156 29988 16158
rect 34300 16156 34356 16212
rect 27468 14642 27524 14644
rect 27468 14590 27470 14642
rect 27470 14590 27522 14642
rect 27522 14590 27524 14642
rect 27468 14588 27524 14590
rect 27580 14306 27636 14308
rect 27580 14254 27582 14306
rect 27582 14254 27634 14306
rect 27634 14254 27636 14306
rect 27580 14252 27636 14254
rect 27132 13746 27188 13748
rect 27132 13694 27134 13746
rect 27134 13694 27186 13746
rect 27186 13694 27188 13746
rect 27132 13692 27188 13694
rect 27020 13468 27076 13524
rect 27468 13468 27524 13524
rect 27244 13020 27300 13076
rect 26908 12012 26964 12068
rect 27020 12124 27076 12180
rect 26796 11900 26852 11956
rect 26012 9772 26068 9828
rect 26012 8988 26068 9044
rect 25676 7532 25732 7588
rect 25788 7420 25844 7476
rect 25564 6748 25620 6804
rect 25676 6524 25732 6580
rect 25676 6076 25732 6132
rect 24556 5292 24612 5348
rect 24780 5628 24836 5684
rect 24668 5234 24724 5236
rect 24668 5182 24670 5234
rect 24670 5182 24722 5234
rect 24722 5182 24724 5234
rect 24668 5180 24724 5182
rect 25900 6300 25956 6356
rect 25788 5068 25844 5124
rect 24892 3836 24948 3892
rect 25340 3612 25396 3668
rect 23996 3388 24052 3444
rect 25452 3442 25508 3444
rect 25452 3390 25454 3442
rect 25454 3390 25506 3442
rect 25506 3390 25508 3442
rect 25452 3388 25508 3390
rect 26236 10108 26292 10164
rect 26684 11452 26740 11508
rect 26572 11170 26628 11172
rect 26572 11118 26574 11170
rect 26574 11118 26626 11170
rect 26626 11118 26628 11170
rect 26572 11116 26628 11118
rect 26796 10498 26852 10500
rect 26796 10446 26798 10498
rect 26798 10446 26850 10498
rect 26850 10446 26852 10498
rect 26796 10444 26852 10446
rect 26684 10220 26740 10276
rect 26460 9772 26516 9828
rect 26348 9436 26404 9492
rect 26124 8204 26180 8260
rect 26236 8876 26292 8932
rect 26236 7308 26292 7364
rect 26236 6636 26292 6692
rect 26460 8204 26516 8260
rect 26460 7532 26516 7588
rect 26796 7420 26852 7476
rect 26684 7362 26740 7364
rect 26684 7310 26686 7362
rect 26686 7310 26738 7362
rect 26738 7310 26740 7362
rect 26684 7308 26740 7310
rect 26572 7084 26628 7140
rect 26796 6972 26852 7028
rect 26460 5292 26516 5348
rect 27244 11788 27300 11844
rect 27132 8428 27188 8484
rect 27020 7868 27076 7924
rect 27132 7196 27188 7252
rect 26684 4956 26740 5012
rect 25788 2716 25844 2772
rect 27468 12850 27524 12852
rect 27468 12798 27470 12850
rect 27470 12798 27522 12850
rect 27522 12798 27524 12850
rect 27468 12796 27524 12798
rect 27468 12290 27524 12292
rect 27468 12238 27470 12290
rect 27470 12238 27522 12290
rect 27522 12238 27524 12290
rect 27468 12236 27524 12238
rect 27692 12796 27748 12852
rect 28252 15372 28308 15428
rect 28028 15314 28084 15316
rect 28028 15262 28030 15314
rect 28030 15262 28082 15314
rect 28082 15262 28084 15314
rect 28028 15260 28084 15262
rect 28028 14642 28084 14644
rect 28028 14590 28030 14642
rect 28030 14590 28082 14642
rect 28082 14590 28084 14642
rect 28028 14588 28084 14590
rect 28140 13970 28196 13972
rect 28140 13918 28142 13970
rect 28142 13918 28194 13970
rect 28194 13918 28196 13970
rect 28140 13916 28196 13918
rect 28140 13244 28196 13300
rect 27916 12908 27972 12964
rect 28476 13244 28532 13300
rect 30716 15538 30772 15540
rect 30716 15486 30718 15538
rect 30718 15486 30770 15538
rect 30770 15486 30772 15538
rect 30716 15484 30772 15486
rect 30044 15372 30100 15428
rect 29820 15314 29876 15316
rect 29820 15262 29822 15314
rect 29822 15262 29874 15314
rect 29874 15262 29876 15314
rect 29820 15260 29876 15262
rect 28812 14252 28868 14308
rect 28924 15148 28980 15204
rect 28812 13692 28868 13748
rect 29036 13916 29092 13972
rect 29372 13634 29428 13636
rect 29372 13582 29374 13634
rect 29374 13582 29426 13634
rect 29426 13582 29428 13634
rect 29372 13580 29428 13582
rect 29484 14252 29540 14308
rect 27804 11900 27860 11956
rect 27356 11340 27412 11396
rect 27356 11170 27412 11172
rect 27356 11118 27358 11170
rect 27358 11118 27410 11170
rect 27410 11118 27412 11170
rect 27356 11116 27412 11118
rect 27468 11004 27524 11060
rect 27468 10668 27524 10724
rect 27356 10444 27412 10500
rect 27580 9996 27636 10052
rect 27468 9938 27524 9940
rect 27468 9886 27470 9938
rect 27470 9886 27522 9938
rect 27522 9886 27524 9938
rect 27468 9884 27524 9886
rect 27804 10050 27860 10052
rect 27804 9998 27806 10050
rect 27806 9998 27858 10050
rect 27858 9998 27860 10050
rect 27804 9996 27860 9998
rect 27692 9324 27748 9380
rect 27692 9100 27748 9156
rect 27580 7698 27636 7700
rect 27580 7646 27582 7698
rect 27582 7646 27634 7698
rect 27634 7646 27636 7698
rect 27580 7644 27636 7646
rect 27804 8930 27860 8932
rect 27804 8878 27806 8930
rect 27806 8878 27858 8930
rect 27858 8878 27860 8930
rect 27804 8876 27860 8878
rect 27804 8204 27860 8260
rect 27692 6412 27748 6468
rect 28364 12460 28420 12516
rect 28812 12460 28868 12516
rect 28812 12236 28868 12292
rect 28364 12012 28420 12068
rect 28252 11900 28308 11956
rect 28700 11564 28756 11620
rect 28588 11452 28644 11508
rect 28588 10780 28644 10836
rect 29372 11900 29428 11956
rect 28476 9938 28532 9940
rect 28476 9886 28478 9938
rect 28478 9886 28530 9938
rect 28530 9886 28532 9938
rect 28476 9884 28532 9886
rect 29260 10668 29316 10724
rect 28588 9042 28644 9044
rect 28588 8990 28590 9042
rect 28590 8990 28642 9042
rect 28642 8990 28644 9042
rect 28588 8988 28644 8990
rect 28252 8204 28308 8260
rect 28588 8316 28644 8372
rect 28252 6748 28308 6804
rect 28476 7474 28532 7476
rect 28476 7422 28478 7474
rect 28478 7422 28530 7474
rect 28530 7422 28532 7474
rect 28476 7420 28532 7422
rect 28588 6018 28644 6020
rect 28588 5966 28590 6018
rect 28590 5966 28642 6018
rect 28642 5966 28644 6018
rect 28588 5964 28644 5966
rect 27804 5180 27860 5236
rect 27468 5010 27524 5012
rect 27468 4958 27470 5010
rect 27470 4958 27522 5010
rect 27522 4958 27524 5010
rect 27468 4956 27524 4958
rect 28700 5068 28756 5124
rect 28476 4508 28532 4564
rect 28924 7084 28980 7140
rect 28924 6188 28980 6244
rect 29148 8764 29204 8820
rect 29260 6972 29316 7028
rect 29932 14306 29988 14308
rect 29932 14254 29934 14306
rect 29934 14254 29986 14306
rect 29986 14254 29988 14306
rect 29932 14252 29988 14254
rect 29820 13746 29876 13748
rect 29820 13694 29822 13746
rect 29822 13694 29874 13746
rect 29874 13694 29876 13746
rect 29820 13692 29876 13694
rect 29596 11564 29652 11620
rect 29484 11004 29540 11060
rect 29484 10108 29540 10164
rect 29036 5964 29092 6020
rect 29372 6130 29428 6132
rect 29372 6078 29374 6130
rect 29374 6078 29426 6130
rect 29426 6078 29428 6130
rect 29372 6076 29428 6078
rect 29036 5068 29092 5124
rect 28812 4284 28868 4340
rect 28588 4226 28644 4228
rect 28588 4174 28590 4226
rect 28590 4174 28642 4226
rect 28642 4174 28644 4226
rect 28588 4172 28644 4174
rect 27804 3666 27860 3668
rect 27804 3614 27806 3666
rect 27806 3614 27858 3666
rect 27858 3614 27860 3666
rect 27804 3612 27860 3614
rect 28028 3612 28084 3668
rect 29820 11564 29876 11620
rect 31164 15426 31220 15428
rect 31164 15374 31166 15426
rect 31166 15374 31218 15426
rect 31218 15374 31220 15426
rect 31164 15372 31220 15374
rect 31948 15260 32004 15316
rect 30380 15202 30436 15204
rect 30380 15150 30382 15202
rect 30382 15150 30434 15202
rect 30434 15150 30436 15202
rect 30380 15148 30436 15150
rect 30268 12850 30324 12852
rect 30268 12798 30270 12850
rect 30270 12798 30322 12850
rect 30322 12798 30324 12850
rect 30268 12796 30324 12798
rect 30268 12572 30324 12628
rect 30156 12178 30212 12180
rect 30156 12126 30158 12178
rect 30158 12126 30210 12178
rect 30210 12126 30212 12178
rect 30156 12124 30212 12126
rect 30940 14306 30996 14308
rect 30940 14254 30942 14306
rect 30942 14254 30994 14306
rect 30994 14254 30996 14306
rect 30940 14252 30996 14254
rect 31612 14306 31668 14308
rect 31612 14254 31614 14306
rect 31614 14254 31666 14306
rect 31666 14254 31668 14306
rect 31612 14252 31668 14254
rect 31164 13634 31220 13636
rect 31164 13582 31166 13634
rect 31166 13582 31218 13634
rect 31218 13582 31220 13634
rect 31164 13580 31220 13582
rect 30716 12684 30772 12740
rect 31276 12796 31332 12852
rect 30604 12012 30660 12068
rect 30380 11788 30436 11844
rect 29932 11394 29988 11396
rect 29932 11342 29934 11394
rect 29934 11342 29986 11394
rect 29986 11342 29988 11394
rect 29932 11340 29988 11342
rect 29820 11116 29876 11172
rect 29708 10332 29764 10388
rect 29596 8988 29652 9044
rect 29708 10108 29764 10164
rect 29596 6972 29652 7028
rect 29820 9212 29876 9268
rect 30268 10668 30324 10724
rect 30380 11116 30436 11172
rect 30044 9826 30100 9828
rect 30044 9774 30046 9826
rect 30046 9774 30098 9826
rect 30098 9774 30100 9826
rect 30044 9772 30100 9774
rect 30380 9436 30436 9492
rect 30044 8316 30100 8372
rect 29820 7196 29876 7252
rect 29932 8204 29988 8260
rect 30268 9154 30324 9156
rect 30268 9102 30270 9154
rect 30270 9102 30322 9154
rect 30322 9102 30324 9154
rect 30268 9100 30324 9102
rect 30268 8930 30324 8932
rect 30268 8878 30270 8930
rect 30270 8878 30322 8930
rect 30322 8878 30324 8930
rect 30268 8876 30324 8878
rect 30940 12066 30996 12068
rect 30940 12014 30942 12066
rect 30942 12014 30994 12066
rect 30994 12014 30996 12066
rect 30940 12012 30996 12014
rect 30828 11954 30884 11956
rect 30828 11902 30830 11954
rect 30830 11902 30882 11954
rect 30882 11902 30884 11954
rect 30828 11900 30884 11902
rect 31052 11452 31108 11508
rect 31052 11282 31108 11284
rect 31052 11230 31054 11282
rect 31054 11230 31106 11282
rect 31106 11230 31108 11282
rect 31052 11228 31108 11230
rect 30716 11116 30772 11172
rect 30492 8204 30548 8260
rect 30604 9996 30660 10052
rect 30268 8034 30324 8036
rect 30268 7982 30270 8034
rect 30270 7982 30322 8034
rect 30322 7982 30324 8034
rect 30268 7980 30324 7982
rect 29932 7644 29988 7700
rect 29820 6466 29876 6468
rect 29820 6414 29822 6466
rect 29822 6414 29874 6466
rect 29874 6414 29876 6466
rect 29820 6412 29876 6414
rect 31052 9772 31108 9828
rect 30940 9436 30996 9492
rect 31164 9714 31220 9716
rect 31164 9662 31166 9714
rect 31166 9662 31218 9714
rect 31218 9662 31220 9714
rect 31164 9660 31220 9662
rect 31724 13804 31780 13860
rect 31948 13916 32004 13972
rect 31500 11954 31556 11956
rect 31500 11902 31502 11954
rect 31502 11902 31554 11954
rect 31554 11902 31556 11954
rect 31500 11900 31556 11902
rect 31388 9772 31444 9828
rect 31500 11452 31556 11508
rect 31052 8876 31108 8932
rect 30940 8818 30996 8820
rect 30940 8766 30942 8818
rect 30942 8766 30994 8818
rect 30994 8766 30996 8818
rect 30940 8764 30996 8766
rect 30604 7980 30660 8036
rect 30492 7308 30548 7364
rect 30604 6690 30660 6692
rect 30604 6638 30606 6690
rect 30606 6638 30658 6690
rect 30658 6638 30660 6690
rect 30604 6636 30660 6638
rect 30492 6578 30548 6580
rect 30492 6526 30494 6578
rect 30494 6526 30546 6578
rect 30546 6526 30548 6578
rect 30492 6524 30548 6526
rect 29596 6188 29652 6244
rect 29932 6018 29988 6020
rect 29932 5966 29934 6018
rect 29934 5966 29986 6018
rect 29986 5966 29988 6018
rect 29932 5964 29988 5966
rect 29820 5906 29876 5908
rect 29820 5854 29822 5906
rect 29822 5854 29874 5906
rect 29874 5854 29876 5906
rect 29820 5852 29876 5854
rect 30380 5906 30436 5908
rect 30380 5854 30382 5906
rect 30382 5854 30434 5906
rect 30434 5854 30436 5906
rect 30380 5852 30436 5854
rect 31836 12012 31892 12068
rect 31724 11676 31780 11732
rect 32620 15202 32676 15204
rect 32620 15150 32622 15202
rect 32622 15150 32674 15202
rect 32674 15150 32676 15202
rect 32620 15148 32676 15150
rect 33740 15148 33796 15204
rect 32844 14476 32900 14532
rect 32396 14306 32452 14308
rect 32396 14254 32398 14306
rect 32398 14254 32450 14306
rect 32450 14254 32452 14306
rect 32396 14252 32452 14254
rect 33292 14418 33348 14420
rect 33292 14366 33294 14418
rect 33294 14366 33346 14418
rect 33346 14366 33348 14418
rect 33292 14364 33348 14366
rect 32172 13970 32228 13972
rect 32172 13918 32174 13970
rect 32174 13918 32226 13970
rect 32226 13918 32228 13970
rect 32172 13916 32228 13918
rect 32284 13804 32340 13860
rect 32172 13132 32228 13188
rect 32172 12236 32228 12292
rect 32620 13634 32676 13636
rect 32620 13582 32622 13634
rect 32622 13582 32674 13634
rect 32674 13582 32676 13634
rect 32620 13580 32676 13582
rect 32396 13132 32452 13188
rect 33404 13580 33460 13636
rect 30828 6972 30884 7028
rect 30940 8092 30996 8148
rect 31388 8258 31444 8260
rect 31388 8206 31390 8258
rect 31390 8206 31442 8258
rect 31442 8206 31444 8258
rect 31388 8204 31444 8206
rect 32060 11564 32116 11620
rect 32060 11170 32116 11172
rect 32060 11118 32062 11170
rect 32062 11118 32114 11170
rect 32114 11118 32116 11170
rect 32060 11116 32116 11118
rect 31724 9996 31780 10052
rect 31836 10444 31892 10500
rect 31724 8988 31780 9044
rect 31836 8930 31892 8932
rect 31836 8878 31838 8930
rect 31838 8878 31890 8930
rect 31890 8878 31892 8930
rect 31836 8876 31892 8878
rect 32060 9436 32116 9492
rect 32956 12460 33012 12516
rect 32732 12290 32788 12292
rect 32732 12238 32734 12290
rect 32734 12238 32786 12290
rect 32786 12238 32788 12290
rect 32732 12236 32788 12238
rect 32844 12178 32900 12180
rect 32844 12126 32846 12178
rect 32846 12126 32898 12178
rect 32898 12126 32900 12178
rect 32844 12124 32900 12126
rect 32396 11676 32452 11732
rect 32620 11452 32676 11508
rect 32396 10498 32452 10500
rect 32396 10446 32398 10498
rect 32398 10446 32450 10498
rect 32450 10446 32452 10498
rect 32396 10444 32452 10446
rect 32620 9324 32676 9380
rect 32508 8988 32564 9044
rect 31948 7868 32004 7924
rect 31276 7362 31332 7364
rect 31276 7310 31278 7362
rect 31278 7310 31330 7362
rect 31330 7310 31332 7362
rect 31276 7308 31332 7310
rect 31052 6076 31108 6132
rect 31164 6860 31220 6916
rect 30716 5234 30772 5236
rect 30716 5182 30718 5234
rect 30718 5182 30770 5234
rect 30770 5182 30772 5234
rect 30716 5180 30772 5182
rect 29932 5122 29988 5124
rect 29932 5070 29934 5122
rect 29934 5070 29986 5122
rect 29986 5070 29988 5122
rect 29932 5068 29988 5070
rect 32508 8316 32564 8372
rect 32844 11170 32900 11172
rect 32844 11118 32846 11170
rect 32846 11118 32898 11170
rect 32898 11118 32900 11170
rect 32844 11116 32900 11118
rect 33292 12124 33348 12180
rect 33180 11394 33236 11396
rect 33180 11342 33182 11394
rect 33182 11342 33234 11394
rect 33234 11342 33236 11394
rect 33180 11340 33236 11342
rect 36540 15372 36596 15428
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 33964 12290 34020 12292
rect 33964 12238 33966 12290
rect 33966 12238 34018 12290
rect 34018 12238 34020 12290
rect 33964 12236 34020 12238
rect 33628 11340 33684 11396
rect 33516 11116 33572 11172
rect 33068 9548 33124 9604
rect 33404 10892 33460 10948
rect 32732 8204 32788 8260
rect 32956 8988 33012 9044
rect 32396 7980 32452 8036
rect 32172 6076 32228 6132
rect 31500 6018 31556 6020
rect 31500 5966 31502 6018
rect 31502 5966 31554 6018
rect 31554 5966 31556 6018
rect 31500 5964 31556 5966
rect 31836 6018 31892 6020
rect 31836 5966 31838 6018
rect 31838 5966 31890 6018
rect 31890 5966 31892 6018
rect 31836 5964 31892 5966
rect 31164 5068 31220 5124
rect 31388 5292 31444 5348
rect 30828 4396 30884 4452
rect 32060 5740 32116 5796
rect 32284 5852 32340 5908
rect 31612 5180 31668 5236
rect 31612 4338 31668 4340
rect 31612 4286 31614 4338
rect 31614 4286 31666 4338
rect 31666 4286 31668 4338
rect 31612 4284 31668 4286
rect 31948 4338 32004 4340
rect 31948 4286 31950 4338
rect 31950 4286 32002 4338
rect 32002 4286 32004 4338
rect 31948 4284 32004 4286
rect 29932 3666 29988 3668
rect 29932 3614 29934 3666
rect 29934 3614 29986 3666
rect 29986 3614 29988 3666
rect 29932 3612 29988 3614
rect 32172 3612 32228 3668
rect 32732 7868 32788 7924
rect 32956 7196 33012 7252
rect 32956 6972 33012 7028
rect 32732 6300 32788 6356
rect 32844 6188 32900 6244
rect 32732 5628 32788 5684
rect 32844 5234 32900 5236
rect 32844 5182 32846 5234
rect 32846 5182 32898 5234
rect 32898 5182 32900 5234
rect 32844 5180 32900 5182
rect 32508 5068 32564 5124
rect 32732 4562 32788 4564
rect 32732 4510 32734 4562
rect 32734 4510 32786 4562
rect 32786 4510 32788 4562
rect 32732 4508 32788 4510
rect 33292 9938 33348 9940
rect 33292 9886 33294 9938
rect 33294 9886 33346 9938
rect 33346 9886 33348 9938
rect 33292 9884 33348 9886
rect 33180 6300 33236 6356
rect 33628 10892 33684 10948
rect 34748 13916 34804 13972
rect 34300 12684 34356 12740
rect 34188 12460 34244 12516
rect 33964 11900 34020 11956
rect 33516 9266 33572 9268
rect 33516 9214 33518 9266
rect 33518 9214 33570 9266
rect 33570 9214 33572 9266
rect 33516 9212 33572 9214
rect 33740 9884 33796 9940
rect 33852 9772 33908 9828
rect 33852 9042 33908 9044
rect 33852 8990 33854 9042
rect 33854 8990 33906 9042
rect 33906 8990 33908 9042
rect 33852 8988 33908 8990
rect 33628 8652 33684 8708
rect 34188 10610 34244 10612
rect 34188 10558 34190 10610
rect 34190 10558 34242 10610
rect 34242 10558 34244 10610
rect 34188 10556 34244 10558
rect 33964 8652 34020 8708
rect 34188 9772 34244 9828
rect 33740 8204 33796 8260
rect 33964 8146 34020 8148
rect 33964 8094 33966 8146
rect 33966 8094 34018 8146
rect 34018 8094 34020 8146
rect 33964 8092 34020 8094
rect 33740 8034 33796 8036
rect 33740 7982 33742 8034
rect 33742 7982 33794 8034
rect 33794 7982 33796 8034
rect 33740 7980 33796 7982
rect 34076 7980 34132 8036
rect 33964 7756 34020 7812
rect 33404 5292 33460 5348
rect 33628 6972 33684 7028
rect 33852 7586 33908 7588
rect 33852 7534 33854 7586
rect 33854 7534 33906 7586
rect 33906 7534 33908 7586
rect 33852 7532 33908 7534
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34748 12572 34804 12628
rect 35532 12850 35588 12852
rect 35532 12798 35534 12850
rect 35534 12798 35586 12850
rect 35586 12798 35588 12850
rect 35532 12796 35588 12798
rect 35084 12738 35140 12740
rect 35084 12686 35086 12738
rect 35086 12686 35138 12738
rect 35138 12686 35140 12738
rect 35084 12684 35140 12686
rect 34972 12460 35028 12516
rect 35084 12236 35140 12292
rect 35532 11954 35588 11956
rect 35532 11902 35534 11954
rect 35534 11902 35586 11954
rect 35586 11902 35588 11954
rect 35532 11900 35588 11902
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34636 11282 34692 11284
rect 34636 11230 34638 11282
rect 34638 11230 34690 11282
rect 34690 11230 34692 11282
rect 34636 11228 34692 11230
rect 34524 10780 34580 10836
rect 34748 9212 34804 9268
rect 34300 8316 34356 8372
rect 34300 7644 34356 7700
rect 34188 6972 34244 7028
rect 34524 8652 34580 8708
rect 34748 8204 34804 8260
rect 34412 6636 34468 6692
rect 33852 6130 33908 6132
rect 33852 6078 33854 6130
rect 33854 6078 33906 6130
rect 33906 6078 33908 6130
rect 33852 6076 33908 6078
rect 33740 5852 33796 5908
rect 34076 5292 34132 5348
rect 33628 5180 33684 5236
rect 33964 5234 34020 5236
rect 33964 5182 33966 5234
rect 33966 5182 34018 5234
rect 34018 5182 34020 5234
rect 33964 5180 34020 5182
rect 33628 4450 33684 4452
rect 33628 4398 33630 4450
rect 33630 4398 33682 4450
rect 33682 4398 33684 4450
rect 33628 4396 33684 4398
rect 33852 4338 33908 4340
rect 33852 4286 33854 4338
rect 33854 4286 33906 4338
rect 33906 4286 33908 4338
rect 33852 4284 33908 4286
rect 34636 6860 34692 6916
rect 34860 7196 34916 7252
rect 35532 10556 35588 10612
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35420 9660 35476 9716
rect 35420 9154 35476 9156
rect 35420 9102 35422 9154
rect 35422 9102 35474 9154
rect 35474 9102 35476 9154
rect 35420 9100 35476 9102
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35868 12460 35924 12516
rect 35756 11676 35812 11732
rect 36428 12738 36484 12740
rect 36428 12686 36430 12738
rect 36430 12686 36482 12738
rect 36482 12686 36484 12738
rect 36428 12684 36484 12686
rect 36652 12684 36708 12740
rect 35644 9660 35700 9716
rect 35644 8988 35700 9044
rect 35084 8204 35140 8260
rect 35532 7868 35588 7924
rect 35532 7586 35588 7588
rect 35532 7534 35534 7586
rect 35534 7534 35586 7586
rect 35586 7534 35588 7586
rect 35532 7532 35588 7534
rect 35084 7196 35140 7252
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 36540 12012 36596 12068
rect 36204 11676 36260 11732
rect 36092 10834 36148 10836
rect 36092 10782 36094 10834
rect 36094 10782 36146 10834
rect 36146 10782 36148 10834
rect 36092 10780 36148 10782
rect 36092 10332 36148 10388
rect 36092 10108 36148 10164
rect 36092 8988 36148 9044
rect 36204 9826 36260 9828
rect 36204 9774 36206 9826
rect 36206 9774 36258 9826
rect 36258 9774 36260 9826
rect 36204 9772 36260 9774
rect 36204 8764 36260 8820
rect 36316 9660 36372 9716
rect 36092 8540 36148 8596
rect 36764 12012 36820 12068
rect 37436 11788 37492 11844
rect 36988 11676 37044 11732
rect 40572 12684 40628 12740
rect 42140 14588 42196 14644
rect 42028 12460 42084 12516
rect 37884 12066 37940 12068
rect 37884 12014 37886 12066
rect 37886 12014 37938 12066
rect 37938 12014 37940 12066
rect 37884 12012 37940 12014
rect 37772 11676 37828 11732
rect 37660 11394 37716 11396
rect 37660 11342 37662 11394
rect 37662 11342 37714 11394
rect 37714 11342 37716 11394
rect 37660 11340 37716 11342
rect 37548 11282 37604 11284
rect 37548 11230 37550 11282
rect 37550 11230 37602 11282
rect 37602 11230 37604 11282
rect 37548 11228 37604 11230
rect 36876 10722 36932 10724
rect 36876 10670 36878 10722
rect 36878 10670 36930 10722
rect 36930 10670 36932 10722
rect 36876 10668 36932 10670
rect 36316 8034 36372 8036
rect 36316 7982 36318 8034
rect 36318 7982 36370 8034
rect 36370 7982 36372 8034
rect 36316 7980 36372 7982
rect 36204 7868 36260 7924
rect 35980 6690 36036 6692
rect 35980 6638 35982 6690
rect 35982 6638 36034 6690
rect 36034 6638 36036 6690
rect 35980 6636 36036 6638
rect 35868 5964 35924 6020
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35980 5346 36036 5348
rect 35980 5294 35982 5346
rect 35982 5294 36034 5346
rect 36034 5294 36036 5346
rect 35980 5292 36036 5294
rect 35420 5068 35476 5124
rect 35084 5010 35140 5012
rect 35084 4958 35086 5010
rect 35086 4958 35138 5010
rect 35138 4958 35140 5010
rect 35084 4956 35140 4958
rect 36428 7644 36484 7700
rect 36316 7196 36372 7252
rect 36988 10108 37044 10164
rect 37996 11788 38052 11844
rect 37772 10444 37828 10500
rect 38220 10834 38276 10836
rect 38220 10782 38222 10834
rect 38222 10782 38274 10834
rect 38274 10782 38276 10834
rect 38220 10780 38276 10782
rect 37996 10610 38052 10612
rect 37996 10558 37998 10610
rect 37998 10558 38050 10610
rect 38050 10558 38052 10610
rect 37996 10556 38052 10558
rect 37436 10108 37492 10164
rect 37660 9938 37716 9940
rect 37660 9886 37662 9938
rect 37662 9886 37714 9938
rect 37714 9886 37716 9938
rect 37660 9884 37716 9886
rect 37436 9324 37492 9380
rect 38108 9826 38164 9828
rect 38108 9774 38110 9826
rect 38110 9774 38162 9826
rect 38162 9774 38164 9826
rect 38108 9772 38164 9774
rect 38220 9660 38276 9716
rect 37548 9100 37604 9156
rect 38220 9324 38276 9380
rect 38668 11394 38724 11396
rect 38668 11342 38670 11394
rect 38670 11342 38722 11394
rect 38722 11342 38724 11394
rect 38668 11340 38724 11342
rect 38556 10556 38612 10612
rect 38780 9996 38836 10052
rect 39004 11394 39060 11396
rect 39004 11342 39006 11394
rect 39006 11342 39058 11394
rect 39058 11342 39060 11394
rect 39004 11340 39060 11342
rect 39228 10780 39284 10836
rect 39676 11340 39732 11396
rect 39564 10780 39620 10836
rect 39004 10556 39060 10612
rect 38668 9938 38724 9940
rect 38668 9886 38670 9938
rect 38670 9886 38722 9938
rect 38722 9886 38724 9938
rect 38668 9884 38724 9886
rect 39116 10668 39172 10724
rect 38444 9772 38500 9828
rect 38780 9714 38836 9716
rect 38780 9662 38782 9714
rect 38782 9662 38834 9714
rect 38834 9662 38836 9714
rect 38780 9660 38836 9662
rect 38556 9548 38612 9604
rect 38444 9042 38500 9044
rect 38444 8990 38446 9042
rect 38446 8990 38498 9042
rect 38498 8990 38500 9042
rect 38444 8988 38500 8990
rect 37548 8930 37604 8932
rect 37548 8878 37550 8930
rect 37550 8878 37602 8930
rect 37602 8878 37604 8930
rect 37548 8876 37604 8878
rect 37996 8540 38052 8596
rect 37660 7532 37716 7588
rect 36876 7308 36932 7364
rect 37660 7362 37716 7364
rect 37660 7310 37662 7362
rect 37662 7310 37714 7362
rect 37714 7310 37716 7362
rect 37660 7308 37716 7310
rect 36652 6860 36708 6916
rect 36764 6802 36820 6804
rect 36764 6750 36766 6802
rect 36766 6750 36818 6802
rect 36818 6750 36820 6802
rect 36764 6748 36820 6750
rect 37884 7420 37940 7476
rect 39004 9714 39060 9716
rect 39004 9662 39006 9714
rect 39006 9662 39058 9714
rect 39058 9662 39060 9714
rect 39004 9660 39060 9662
rect 40236 10780 40292 10836
rect 39788 10556 39844 10612
rect 40124 10610 40180 10612
rect 40124 10558 40126 10610
rect 40126 10558 40178 10610
rect 40178 10558 40180 10610
rect 40124 10556 40180 10558
rect 39676 10332 39732 10388
rect 39228 10220 39284 10276
rect 39788 10220 39844 10276
rect 39564 9714 39620 9716
rect 39564 9662 39566 9714
rect 39566 9662 39618 9714
rect 39618 9662 39620 9714
rect 39564 9660 39620 9662
rect 40124 9826 40180 9828
rect 40124 9774 40126 9826
rect 40126 9774 40178 9826
rect 40178 9774 40180 9826
rect 40124 9772 40180 9774
rect 39676 8988 39732 9044
rect 40012 8988 40068 9044
rect 39004 8876 39060 8932
rect 38668 8764 38724 8820
rect 39340 8540 39396 8596
rect 39564 8370 39620 8372
rect 39564 8318 39566 8370
rect 39566 8318 39618 8370
rect 39618 8318 39620 8370
rect 39564 8316 39620 8318
rect 39228 8258 39284 8260
rect 39228 8206 39230 8258
rect 39230 8206 39282 8258
rect 39282 8206 39284 8258
rect 39228 8204 39284 8206
rect 38220 7980 38276 8036
rect 38332 7698 38388 7700
rect 38332 7646 38334 7698
rect 38334 7646 38386 7698
rect 38386 7646 38388 7698
rect 38332 7644 38388 7646
rect 37660 6076 37716 6132
rect 37548 5964 37604 6020
rect 37436 5852 37492 5908
rect 36092 4172 36148 4228
rect 33852 3666 33908 3668
rect 33852 3614 33854 3666
rect 33854 3614 33906 3666
rect 33906 3614 33908 3666
rect 33852 3612 33908 3614
rect 33404 3500 33460 3556
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35644 3500 35700 3556
rect 34748 3388 34804 3444
rect 38108 6076 38164 6132
rect 38332 5628 38388 5684
rect 37884 5292 37940 5348
rect 38556 7420 38612 7476
rect 38444 5292 38500 5348
rect 37884 5068 37940 5124
rect 38220 4226 38276 4228
rect 38220 4174 38222 4226
rect 38222 4174 38274 4226
rect 38274 4174 38276 4226
rect 38220 4172 38276 4174
rect 38332 4060 38388 4116
rect 37212 3442 37268 3444
rect 37212 3390 37214 3442
rect 37214 3390 37266 3442
rect 37266 3390 37268 3442
rect 37212 3388 37268 3390
rect 37436 3388 37492 3444
rect 39340 5906 39396 5908
rect 39340 5854 39342 5906
rect 39342 5854 39394 5906
rect 39394 5854 39396 5906
rect 39340 5852 39396 5854
rect 39788 7868 39844 7924
rect 39788 7532 39844 7588
rect 39676 7308 39732 7364
rect 39564 6018 39620 6020
rect 39564 5966 39566 6018
rect 39566 5966 39618 6018
rect 39618 5966 39620 6018
rect 39564 5964 39620 5966
rect 40124 8370 40180 8372
rect 40124 8318 40126 8370
rect 40126 8318 40178 8370
rect 40178 8318 40180 8370
rect 40124 8316 40180 8318
rect 40572 10834 40628 10836
rect 40572 10782 40574 10834
rect 40574 10782 40626 10834
rect 40626 10782 40628 10834
rect 40572 10780 40628 10782
rect 41356 10556 41412 10612
rect 40572 9996 40628 10052
rect 41020 9826 41076 9828
rect 41020 9774 41022 9826
rect 41022 9774 41074 9826
rect 41074 9774 41076 9826
rect 41020 9772 41076 9774
rect 40460 8428 40516 8484
rect 40684 8428 40740 8484
rect 41244 8316 41300 8372
rect 40684 8034 40740 8036
rect 40684 7982 40686 8034
rect 40686 7982 40738 8034
rect 40738 7982 40740 8034
rect 40684 7980 40740 7982
rect 40348 7868 40404 7924
rect 40236 7644 40292 7700
rect 40124 6690 40180 6692
rect 40124 6638 40126 6690
rect 40126 6638 40178 6690
rect 40178 6638 40180 6690
rect 40124 6636 40180 6638
rect 40796 7250 40852 7252
rect 40796 7198 40798 7250
rect 40798 7198 40850 7250
rect 40850 7198 40852 7250
rect 40796 7196 40852 7198
rect 41132 8146 41188 8148
rect 41132 8094 41134 8146
rect 41134 8094 41186 8146
rect 41186 8094 41188 8146
rect 41132 8092 41188 8094
rect 40348 5964 40404 6020
rect 40908 6076 40964 6132
rect 41020 7980 41076 8036
rect 41020 6748 41076 6804
rect 39452 5068 39508 5124
rect 40124 5180 40180 5236
rect 40012 4562 40068 4564
rect 40012 4510 40014 4562
rect 40014 4510 40066 4562
rect 40066 4510 40068 4562
rect 40012 4508 40068 4510
rect 39340 4396 39396 4452
rect 39900 4114 39956 4116
rect 39900 4062 39902 4114
rect 39902 4062 39954 4114
rect 39954 4062 39956 4114
rect 39900 4060 39956 4062
rect 39228 3836 39284 3892
rect 40684 5122 40740 5124
rect 40684 5070 40686 5122
rect 40686 5070 40738 5122
rect 40738 5070 40740 5122
rect 40684 5068 40740 5070
rect 41804 10444 41860 10500
rect 41468 8316 41524 8372
rect 41580 10108 41636 10164
rect 41916 10220 41972 10276
rect 41916 9548 41972 9604
rect 41692 7362 41748 7364
rect 41692 7310 41694 7362
rect 41694 7310 41746 7362
rect 41746 7310 41748 7362
rect 41692 7308 41748 7310
rect 41580 7250 41636 7252
rect 41580 7198 41582 7250
rect 41582 7198 41634 7250
rect 41634 7198 41636 7250
rect 41580 7196 41636 7198
rect 41692 6636 41748 6692
rect 42028 8034 42084 8036
rect 42028 7982 42030 8034
rect 42030 7982 42082 8034
rect 42082 7982 42084 8034
rect 42028 7980 42084 7982
rect 41916 6188 41972 6244
rect 42028 6466 42084 6468
rect 42028 6414 42030 6466
rect 42030 6414 42082 6466
rect 42082 6414 42084 6466
rect 42028 6412 42084 6414
rect 41804 6130 41860 6132
rect 41804 6078 41806 6130
rect 41806 6078 41858 6130
rect 41858 6078 41860 6130
rect 41804 6076 41860 6078
rect 41804 5292 41860 5348
rect 41356 5234 41412 5236
rect 41356 5182 41358 5234
rect 41358 5182 41410 5234
rect 41410 5182 41412 5234
rect 41356 5180 41412 5182
rect 41244 4508 41300 4564
rect 41692 4508 41748 4564
rect 41580 4450 41636 4452
rect 41580 4398 41582 4450
rect 41582 4398 41634 4450
rect 41634 4398 41636 4450
rect 41580 4396 41636 4398
rect 39116 3612 39172 3668
rect 40908 3724 40964 3780
rect 39004 3442 39060 3444
rect 39004 3390 39006 3442
rect 39006 3390 39058 3442
rect 39058 3390 39060 3442
rect 39004 3388 39060 3390
rect 41468 3612 41524 3668
rect 40124 3554 40180 3556
rect 40124 3502 40126 3554
rect 40126 3502 40178 3554
rect 40178 3502 40180 3554
rect 40124 3500 40180 3502
rect 41580 3500 41636 3556
rect 41916 4956 41972 5012
rect 42476 19852 42532 19908
rect 42364 19740 42420 19796
rect 42364 6748 42420 6804
rect 42140 4620 42196 4676
rect 42364 2940 42420 2996
rect 42588 3276 42644 3332
rect 42476 2828 42532 2884
rect 42812 12460 42868 12516
rect 42812 6412 42868 6468
rect 42924 6748 42980 6804
rect 42700 2604 42756 2660
rect 42812 3836 42868 3892
rect 42924 2492 42980 2548
<< metal3 >>
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 0 33012 800 33040
rect 0 32956 980 33012
rect 0 32928 800 32956
rect 924 32676 980 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 700 32620 980 32676
rect 700 32340 756 32620
rect 700 32284 15932 32340
rect 15988 32284 15998 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 2482 25452 2492 25508
rect 2548 25452 6860 25508
rect 6916 25452 6926 25508
rect 1698 25340 1708 25396
rect 1764 25340 13468 25396
rect 13524 25340 13534 25396
rect 1474 25228 1484 25284
rect 1540 25228 2940 25284
rect 2996 25228 3006 25284
rect 9538 25228 9548 25284
rect 9604 25228 20972 25284
rect 21028 25228 21038 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 2258 24668 2268 24724
rect 2324 24668 6860 24724
rect 6916 24668 6926 24724
rect 2706 24556 2716 24612
rect 2772 24556 4956 24612
rect 5012 24556 5022 24612
rect 11078 24556 11116 24612
rect 11172 24556 11182 24612
rect 3826 24444 3836 24500
rect 3892 24444 7644 24500
rect 7700 24444 9548 24500
rect 9604 24444 9614 24500
rect 11218 24332 11228 24388
rect 11284 24332 11564 24388
rect 11620 24332 14476 24388
rect 14532 24332 14542 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 9986 24220 9996 24276
rect 10052 24220 19516 24276
rect 19572 24220 19582 24276
rect 6402 24108 6412 24164
rect 6468 24108 9156 24164
rect 14018 24108 14028 24164
rect 14084 24108 23548 24164
rect 23604 24108 23614 24164
rect 9100 24052 9156 24108
rect 6178 23996 6188 24052
rect 6244 23996 8652 24052
rect 8708 23996 8718 24052
rect 9090 23996 9100 24052
rect 9156 23996 10780 24052
rect 10836 23996 12236 24052
rect 12292 23996 12302 24052
rect 13458 23996 13468 24052
rect 13524 23996 15036 24052
rect 15092 23996 19404 24052
rect 19460 23996 19470 24052
rect 3266 23884 3276 23940
rect 3332 23884 5964 23940
rect 6020 23884 6030 23940
rect 8092 23884 11452 23940
rect 11508 23884 11518 23940
rect 13570 23884 13580 23940
rect 13636 23884 42700 23940
rect 42756 23884 42766 23940
rect 8092 23828 8148 23884
rect 1586 23772 1596 23828
rect 1652 23772 3724 23828
rect 3780 23772 3790 23828
rect 5730 23772 5740 23828
rect 5796 23772 8148 23828
rect 8306 23772 8316 23828
rect 8372 23772 17612 23828
rect 17668 23772 17678 23828
rect 1362 23660 1372 23716
rect 1428 23660 1932 23716
rect 1988 23660 1998 23716
rect 4274 23660 4284 23716
rect 4340 23660 4620 23716
rect 4676 23660 4686 23716
rect 4946 23660 4956 23716
rect 5012 23660 12684 23716
rect 12740 23660 12750 23716
rect 1138 23548 1148 23604
rect 1204 23548 3276 23604
rect 3332 23548 3342 23604
rect 3826 23548 3836 23604
rect 3892 23548 6860 23604
rect 6916 23548 6926 23604
rect 7830 23548 7868 23604
rect 7924 23548 7934 23604
rect 9650 23548 9660 23604
rect 9716 23548 10892 23604
rect 10948 23548 11676 23604
rect 11732 23548 11742 23604
rect 11890 23548 11900 23604
rect 11956 23548 13804 23604
rect 13860 23548 13870 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 4386 23436 4396 23492
rect 4452 23436 7420 23492
rect 7476 23436 8764 23492
rect 8820 23436 8830 23492
rect 2146 23324 2156 23380
rect 2212 23324 3052 23380
rect 3108 23324 5740 23380
rect 5796 23324 5806 23380
rect 3332 23212 9716 23268
rect 9874 23212 9884 23268
rect 9940 23212 10668 23268
rect 10724 23212 10734 23268
rect 3332 23156 3388 23212
rect 8204 23156 8260 23212
rect 9660 23156 9716 23212
rect 2706 23100 2716 23156
rect 2772 23100 3388 23156
rect 6290 23100 6300 23156
rect 6356 23100 6860 23156
rect 6916 23100 7420 23156
rect 7476 23100 7486 23156
rect 8194 23100 8204 23156
rect 8260 23100 8270 23156
rect 9660 23100 10220 23156
rect 10276 23100 13020 23156
rect 13076 23100 14028 23156
rect 14084 23100 14094 23156
rect 16818 23100 16828 23156
rect 16884 23100 21308 23156
rect 21364 23100 21374 23156
rect 1782 22988 1820 23044
rect 1876 22988 1886 23044
rect 2566 22988 2604 23044
rect 2660 22988 5404 23044
rect 5460 22988 5470 23044
rect 6402 22988 6412 23044
rect 6468 22988 7868 23044
rect 7924 22988 7934 23044
rect 12674 22988 12684 23044
rect 12740 22988 13804 23044
rect 13860 22988 16940 23044
rect 16996 22988 17006 23044
rect 3154 22876 3164 22932
rect 3220 22876 6020 22932
rect 6514 22876 6524 22932
rect 6580 22876 8092 22932
rect 8148 22876 8540 22932
rect 8596 22876 8606 22932
rect 10658 22876 10668 22932
rect 10724 22876 13468 22932
rect 13524 22876 13534 22932
rect 5964 22820 6020 22876
rect 5964 22764 12236 22820
rect 12292 22764 16492 22820
rect 16548 22764 16828 22820
rect 16884 22764 16894 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 6178 22652 6188 22708
rect 6244 22652 7420 22708
rect 7476 22652 7486 22708
rect 1810 22540 1820 22596
rect 1876 22540 10108 22596
rect 10164 22540 10174 22596
rect 17826 22540 17836 22596
rect 17892 22540 42588 22596
rect 42644 22540 42654 22596
rect 4834 22428 4844 22484
rect 4900 22428 6076 22484
rect 6132 22428 6142 22484
rect 10882 22428 10892 22484
rect 10948 22428 11340 22484
rect 11396 22428 11406 22484
rect 17378 22428 17388 22484
rect 17444 22428 42252 22484
rect 42308 22428 42318 22484
rect 1250 22316 1260 22372
rect 1316 22316 4060 22372
rect 4116 22316 4126 22372
rect 9986 22316 9996 22372
rect 10052 22316 10556 22372
rect 10612 22316 10622 22372
rect 16034 22316 16044 22372
rect 16100 22316 25340 22372
rect 25396 22316 25406 22372
rect 39106 22316 39116 22372
rect 39172 22316 40572 22372
rect 40628 22316 40638 22372
rect 5730 22204 5740 22260
rect 5796 22204 6300 22260
rect 6356 22204 6366 22260
rect 9202 22204 9212 22260
rect 9268 22204 10108 22260
rect 10164 22204 10174 22260
rect 14018 22204 14028 22260
rect 14084 22204 15148 22260
rect 15204 22204 16492 22260
rect 16548 22204 18060 22260
rect 18116 22204 18126 22260
rect 2080 22092 2156 22148
rect 2212 22092 5516 22148
rect 5572 22092 5582 22148
rect 8530 22092 8540 22148
rect 8596 22092 8764 22148
rect 8820 22092 10444 22148
rect 10500 22092 10510 22148
rect 12338 22092 12348 22148
rect 12404 22092 12684 22148
rect 12740 22092 13132 22148
rect 13188 22092 13198 22148
rect 14130 22092 14140 22148
rect 14196 22092 15372 22148
rect 15428 22092 16156 22148
rect 16212 22092 16222 22148
rect 16930 22092 16940 22148
rect 16996 22092 18284 22148
rect 18340 22092 22316 22148
rect 22372 22092 22382 22148
rect 43200 22036 44000 22064
rect 7186 21980 7196 22036
rect 7252 21980 10668 22036
rect 10724 21980 10734 22036
rect 40002 21980 40012 22036
rect 40068 21980 44000 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 43200 21952 44000 21980
rect 6486 21868 6524 21924
rect 6580 21868 6590 21924
rect 6850 21868 6860 21924
rect 6916 21868 7420 21924
rect 7476 21868 9772 21924
rect 9828 21868 11004 21924
rect 11060 21868 11070 21924
rect 12338 21868 12348 21924
rect 12404 21868 12908 21924
rect 12964 21868 14140 21924
rect 14196 21868 14206 21924
rect 15474 21868 15484 21924
rect 15540 21868 15820 21924
rect 15876 21868 15886 21924
rect 16146 21868 16156 21924
rect 16212 21868 18284 21924
rect 18340 21868 18350 21924
rect 1922 21756 1932 21812
rect 1988 21756 3836 21812
rect 3892 21756 3902 21812
rect 4050 21756 4060 21812
rect 4116 21756 4732 21812
rect 4788 21756 4798 21812
rect 5730 21756 5740 21812
rect 5796 21756 9100 21812
rect 9156 21756 9166 21812
rect 10070 21756 10108 21812
rect 10164 21756 10174 21812
rect 10546 21756 10556 21812
rect 10612 21756 11564 21812
rect 11620 21756 11788 21812
rect 11844 21756 11854 21812
rect 17602 21756 17612 21812
rect 17668 21756 20300 21812
rect 20356 21756 20366 21812
rect 5740 21700 5796 21756
rect 4274 21644 4284 21700
rect 4340 21644 4844 21700
rect 4900 21644 5796 21700
rect 9538 21644 9548 21700
rect 9604 21644 10668 21700
rect 10724 21644 10734 21700
rect 14914 21644 14924 21700
rect 14980 21644 16044 21700
rect 16100 21644 16492 21700
rect 16548 21644 16558 21700
rect 3798 21532 3836 21588
rect 3892 21532 3902 21588
rect 5394 21532 5404 21588
rect 5460 21532 8092 21588
rect 8148 21532 14700 21588
rect 14756 21532 16156 21588
rect 16212 21532 16222 21588
rect 3490 21420 3500 21476
rect 3556 21420 5628 21476
rect 5684 21420 5694 21476
rect 7410 21420 7420 21476
rect 7476 21420 7532 21476
rect 7588 21420 7598 21476
rect 12002 21420 12012 21476
rect 12068 21420 15372 21476
rect 15428 21420 15438 21476
rect 18134 21420 18172 21476
rect 18228 21420 18238 21476
rect 18498 21420 18508 21476
rect 18564 21420 18620 21476
rect 18676 21420 18686 21476
rect 18172 21364 18228 21420
rect 6514 21308 6524 21364
rect 6580 21308 18228 21364
rect 8306 21196 8316 21252
rect 8372 21196 14476 21252
rect 14532 21196 14542 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 6626 21084 6636 21140
rect 6692 21084 6748 21140
rect 6804 21084 14308 21140
rect 7522 20972 7532 21028
rect 7588 20972 7644 21028
rect 7700 20972 7710 21028
rect 14252 20916 14308 21084
rect 14466 20972 14476 21028
rect 14532 20972 14924 21028
rect 14980 20972 14990 21028
rect 4946 20860 4956 20916
rect 5012 20860 7084 20916
rect 7140 20860 8988 20916
rect 9044 20860 11564 20916
rect 11620 20860 11900 20916
rect 11956 20860 11966 20916
rect 14252 20860 20524 20916
rect 20580 20860 20590 20916
rect 4722 20748 4732 20804
rect 4788 20748 5516 20804
rect 5572 20748 5582 20804
rect 6626 20748 6636 20804
rect 6692 20748 12124 20804
rect 12180 20748 12908 20804
rect 12964 20748 12974 20804
rect 2034 20636 2044 20692
rect 2100 20636 2604 20692
rect 2660 20636 3500 20692
rect 3556 20636 3566 20692
rect 3938 20636 3948 20692
rect 4004 20636 7756 20692
rect 7812 20636 7980 20692
rect 8036 20636 8428 20692
rect 8484 20636 8494 20692
rect 15092 20636 19628 20692
rect 19684 20636 19694 20692
rect 15092 20580 15148 20636
rect 2930 20524 2940 20580
rect 2996 20524 4620 20580
rect 4676 20524 6300 20580
rect 6356 20524 6366 20580
rect 7634 20524 7644 20580
rect 7700 20524 7980 20580
rect 8036 20524 8046 20580
rect 8530 20524 8540 20580
rect 8596 20524 9100 20580
rect 9156 20524 9324 20580
rect 9380 20524 10220 20580
rect 10276 20524 10286 20580
rect 12422 20524 12460 20580
rect 12516 20524 15148 20580
rect 16258 20524 16268 20580
rect 16324 20524 16940 20580
rect 16996 20524 17006 20580
rect 17910 20524 17948 20580
rect 18004 20524 18014 20580
rect 18722 20524 18732 20580
rect 18788 20524 22540 20580
rect 22596 20524 22606 20580
rect 17948 20468 18004 20524
rect 3602 20412 3612 20468
rect 3668 20412 3948 20468
rect 4004 20412 4014 20468
rect 5954 20412 5964 20468
rect 6020 20412 7196 20468
rect 7252 20412 7262 20468
rect 9874 20412 9884 20468
rect 9940 20412 18004 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 3714 20300 3724 20356
rect 3780 20300 7644 20356
rect 7700 20300 7710 20356
rect 16146 20300 16156 20356
rect 16212 20300 17388 20356
rect 17444 20300 17454 20356
rect 2258 20188 2268 20244
rect 2324 20188 2380 20244
rect 2436 20188 2446 20244
rect 2706 20188 2716 20244
rect 2772 20188 3276 20244
rect 3332 20188 4060 20244
rect 4116 20188 4126 20244
rect 4274 20188 4284 20244
rect 4340 20188 6076 20244
rect 6132 20188 6142 20244
rect 10658 20188 10668 20244
rect 10724 20188 11340 20244
rect 11396 20188 11406 20244
rect 12898 20188 12908 20244
rect 12964 20188 16604 20244
rect 16660 20188 19852 20244
rect 19908 20188 19918 20244
rect 5618 20076 5628 20132
rect 5684 20076 7868 20132
rect 7924 20076 10892 20132
rect 10948 20076 12460 20132
rect 12516 20076 13356 20132
rect 13412 20076 15036 20132
rect 15092 20076 15102 20132
rect 15922 20076 15932 20132
rect 15988 20076 18172 20132
rect 18228 20076 18238 20132
rect 2482 19964 2492 20020
rect 2548 19964 2828 20020
rect 2884 19964 8540 20020
rect 8596 19964 8606 20020
rect 9202 19964 9212 20020
rect 9268 19964 9436 20020
rect 9492 19964 10444 20020
rect 10500 19964 12348 20020
rect 12404 19964 12414 20020
rect 10892 19908 10948 19964
rect 5058 19852 5068 19908
rect 5124 19852 6412 19908
rect 6468 19852 7196 19908
rect 7252 19852 7262 19908
rect 10882 19852 10892 19908
rect 10948 19852 10958 19908
rect 12002 19852 12012 19908
rect 12068 19852 14028 19908
rect 14084 19852 14094 19908
rect 16678 19852 16716 19908
rect 16772 19852 16782 19908
rect 17602 19852 17612 19908
rect 17668 19852 19292 19908
rect 19348 19852 19358 19908
rect 20066 19852 20076 19908
rect 20132 19852 42476 19908
rect 42532 19852 42542 19908
rect 4050 19740 4060 19796
rect 4116 19740 6748 19796
rect 6804 19740 7084 19796
rect 7140 19740 7150 19796
rect 8866 19740 8876 19796
rect 8932 19740 9436 19796
rect 9492 19740 9502 19796
rect 9650 19740 9660 19796
rect 9716 19740 16940 19796
rect 16996 19740 17006 19796
rect 21410 19740 21420 19796
rect 21476 19740 42364 19796
rect 42420 19740 42430 19796
rect 5954 19628 5964 19684
rect 6020 19628 22428 19684
rect 22484 19628 22494 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 6514 19516 6524 19572
rect 6580 19516 6860 19572
rect 6916 19516 6926 19572
rect 15474 19516 15484 19572
rect 15540 19516 18620 19572
rect 18676 19516 18686 19572
rect 1922 19404 1932 19460
rect 1988 19404 2156 19460
rect 2212 19404 3500 19460
rect 3556 19404 3566 19460
rect 5058 19404 5068 19460
rect 5124 19404 5180 19460
rect 5236 19404 5246 19460
rect 7084 19404 8092 19460
rect 8148 19404 8316 19460
rect 8372 19404 8382 19460
rect 8754 19404 8764 19460
rect 8820 19404 9212 19460
rect 9268 19404 9278 19460
rect 11666 19404 11676 19460
rect 11732 19404 12572 19460
rect 12628 19404 13580 19460
rect 13636 19404 14252 19460
rect 14308 19404 14318 19460
rect 7084 19348 7140 19404
rect 7074 19292 7084 19348
rect 7140 19292 7150 19348
rect 8194 19292 8204 19348
rect 8260 19292 9100 19348
rect 9156 19292 17836 19348
rect 17892 19292 17902 19348
rect 18050 19292 18060 19348
rect 18116 19292 19404 19348
rect 19460 19292 19470 19348
rect 20290 19292 20300 19348
rect 20356 19292 23548 19348
rect 23604 19292 23614 19348
rect 6514 19180 6524 19236
rect 6580 19180 6636 19236
rect 6692 19180 6702 19236
rect 9874 19180 9884 19236
rect 9940 19180 10444 19236
rect 10500 19180 16716 19236
rect 16772 19180 16782 19236
rect 2258 19068 2268 19124
rect 2324 19068 2492 19124
rect 2548 19068 2558 19124
rect 7634 19068 7644 19124
rect 7700 19068 8092 19124
rect 8148 19068 10108 19124
rect 10164 19068 10668 19124
rect 10724 19068 10734 19124
rect 14914 19068 14924 19124
rect 14980 19068 18508 19124
rect 18564 19068 18956 19124
rect 19012 19068 19022 19124
rect 2146 18956 2156 19012
rect 2212 18956 2716 19012
rect 2772 18956 3612 19012
rect 3668 18956 3678 19012
rect 8950 18956 8988 19012
rect 9044 18956 9054 19012
rect 12002 18956 12012 19012
rect 12068 18956 12684 19012
rect 12740 18956 12750 19012
rect 14130 18956 14140 19012
rect 14196 18956 14588 19012
rect 14644 18956 14924 19012
rect 14980 18956 14990 19012
rect 16034 18956 16044 19012
rect 16100 18956 16380 19012
rect 16436 18956 17388 19012
rect 17444 18956 17454 19012
rect 19842 18956 19852 19012
rect 19908 18956 20188 19012
rect 20244 18956 20254 19012
rect 4610 18844 4620 18900
rect 4676 18844 5068 18900
rect 5124 18844 5134 18900
rect 14140 18788 14196 18956
rect 16818 18844 16828 18900
rect 16884 18844 16940 18900
rect 16996 18844 17006 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 5058 18732 5068 18788
rect 5124 18732 6524 18788
rect 6580 18732 6590 18788
rect 11778 18732 11788 18788
rect 11844 18732 12684 18788
rect 12740 18732 14196 18788
rect 6626 18620 6636 18676
rect 6692 18620 7868 18676
rect 7924 18620 8092 18676
rect 8148 18620 8158 18676
rect 8306 18620 8316 18676
rect 8372 18620 9884 18676
rect 9940 18620 9950 18676
rect 10434 18620 10444 18676
rect 10500 18620 10892 18676
rect 10948 18620 10958 18676
rect 11218 18620 11228 18676
rect 11284 18620 14084 18676
rect 14242 18620 14252 18676
rect 14308 18620 15708 18676
rect 15764 18620 18060 18676
rect 18116 18620 18126 18676
rect 11228 18564 11284 18620
rect 14028 18564 14084 18620
rect 4918 18508 4956 18564
rect 5012 18508 5022 18564
rect 6402 18508 6412 18564
rect 6468 18508 7532 18564
rect 7588 18508 8148 18564
rect 8530 18508 8540 18564
rect 8596 18508 9772 18564
rect 9828 18508 9838 18564
rect 10994 18508 11004 18564
rect 11060 18508 11284 18564
rect 11890 18508 11900 18564
rect 11956 18508 12236 18564
rect 12292 18508 12302 18564
rect 12898 18508 12908 18564
rect 12964 18508 13244 18564
rect 13300 18508 13310 18564
rect 14018 18508 14028 18564
rect 14084 18508 14700 18564
rect 14756 18508 15036 18564
rect 15092 18508 15102 18564
rect 17042 18508 17052 18564
rect 17108 18508 17612 18564
rect 17668 18508 17678 18564
rect 19170 18508 19180 18564
rect 19236 18508 22876 18564
rect 22932 18508 22942 18564
rect 8092 18452 8148 18508
rect 1810 18396 1820 18452
rect 1876 18396 1932 18452
rect 1988 18396 1998 18452
rect 3378 18396 3388 18452
rect 3444 18396 5964 18452
rect 6020 18396 6356 18452
rect 6486 18396 6524 18452
rect 6580 18396 6590 18452
rect 8092 18396 8540 18452
rect 8596 18396 8606 18452
rect 9426 18396 9436 18452
rect 9492 18396 13468 18452
rect 13524 18396 14588 18452
rect 14644 18396 14654 18452
rect 18162 18396 18172 18452
rect 18228 18396 18508 18452
rect 18564 18396 18574 18452
rect 19058 18396 19068 18452
rect 19124 18396 22876 18452
rect 22932 18396 22942 18452
rect 6300 18340 6356 18396
rect 1698 18284 1708 18340
rect 1764 18284 2044 18340
rect 2100 18284 2156 18340
rect 2212 18284 2222 18340
rect 3154 18284 3164 18340
rect 3220 18284 4284 18340
rect 4340 18284 4350 18340
rect 4834 18284 4844 18340
rect 4900 18284 5292 18340
rect 5348 18284 5358 18340
rect 6300 18284 6412 18340
rect 6468 18284 6478 18340
rect 7522 18284 7532 18340
rect 7588 18284 11564 18340
rect 11620 18284 11630 18340
rect 12786 18284 12796 18340
rect 12852 18284 12908 18340
rect 12964 18284 12974 18340
rect 14802 18284 14812 18340
rect 14868 18284 15596 18340
rect 15652 18284 15662 18340
rect 19170 18284 19180 18340
rect 19236 18284 20188 18340
rect 20244 18284 20254 18340
rect 21074 18284 21084 18340
rect 21140 18284 22652 18340
rect 22708 18284 22718 18340
rect 4844 18228 4900 18284
rect 2370 18172 2380 18228
rect 2436 18172 4900 18228
rect 5292 18228 5348 18284
rect 5292 18172 5404 18228
rect 5460 18172 7532 18228
rect 7588 18172 7980 18228
rect 8036 18172 8046 18228
rect 9846 18172 9884 18228
rect 9940 18172 9950 18228
rect 10882 18172 10892 18228
rect 10948 18172 11452 18228
rect 11508 18172 11518 18228
rect 12338 18172 12348 18228
rect 12404 18172 12796 18228
rect 12852 18172 15820 18228
rect 15876 18172 17388 18228
rect 17444 18172 17454 18228
rect 20178 18172 20188 18228
rect 20244 18172 25228 18228
rect 25284 18172 25294 18228
rect 3714 18060 3724 18116
rect 3780 18060 3948 18116
rect 4004 18060 4014 18116
rect 6402 18060 6412 18116
rect 6468 18060 6636 18116
rect 6692 18060 21868 18116
rect 21924 18060 21934 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5842 17948 5852 18004
rect 5908 17948 7196 18004
rect 7252 17948 9660 18004
rect 9716 17948 9726 18004
rect 13010 17948 13020 18004
rect 13076 17948 15148 18004
rect 15204 17948 15708 18004
rect 15764 17948 16156 18004
rect 16212 17948 16222 18004
rect 3042 17836 3052 17892
rect 3108 17836 6300 17892
rect 6356 17836 6366 17892
rect 8194 17836 8204 17892
rect 8260 17836 8428 17892
rect 8484 17836 8494 17892
rect 15362 17836 15372 17892
rect 15428 17836 16492 17892
rect 16548 17836 16828 17892
rect 16884 17836 16894 17892
rect 19282 17836 19292 17892
rect 19348 17836 20300 17892
rect 20356 17836 20860 17892
rect 20916 17836 20926 17892
rect 2706 17724 2716 17780
rect 2772 17724 7420 17780
rect 7476 17724 7486 17780
rect 13346 17724 13356 17780
rect 13412 17724 14140 17780
rect 14196 17724 14206 17780
rect 23538 17724 23548 17780
rect 23604 17724 23884 17780
rect 23940 17724 23950 17780
rect 2594 17612 2604 17668
rect 2660 17612 3276 17668
rect 3332 17612 4396 17668
rect 4452 17612 4462 17668
rect 5618 17612 5628 17668
rect 5684 17612 6356 17668
rect 6514 17612 6524 17668
rect 6580 17612 7196 17668
rect 7252 17612 7262 17668
rect 7494 17612 7532 17668
rect 7588 17612 7598 17668
rect 8194 17612 8204 17668
rect 8260 17612 10332 17668
rect 10388 17612 10398 17668
rect 12114 17612 12124 17668
rect 12180 17612 12460 17668
rect 12516 17612 12684 17668
rect 12740 17612 12750 17668
rect 14466 17612 14476 17668
rect 14532 17612 15372 17668
rect 15428 17612 15438 17668
rect 20178 17612 20188 17668
rect 20244 17612 21532 17668
rect 21588 17612 21598 17668
rect 6300 17556 6356 17612
rect 2706 17500 2716 17556
rect 2772 17500 2828 17556
rect 2884 17500 6076 17556
rect 6132 17500 6142 17556
rect 6300 17500 8540 17556
rect 8596 17500 9884 17556
rect 9940 17500 9950 17556
rect 11218 17500 11228 17556
rect 11284 17500 11676 17556
rect 11732 17500 11742 17556
rect 12898 17500 12908 17556
rect 12964 17500 19068 17556
rect 19124 17500 19134 17556
rect 3042 17388 3052 17444
rect 3108 17388 4172 17444
rect 4228 17388 4844 17444
rect 4900 17388 4910 17444
rect 5058 17388 5068 17444
rect 5124 17388 5292 17444
rect 5348 17388 5684 17444
rect 5842 17388 5852 17444
rect 5908 17388 7420 17444
rect 7476 17388 7486 17444
rect 9174 17388 9212 17444
rect 9268 17388 9278 17444
rect 9650 17388 9660 17444
rect 9716 17388 12796 17444
rect 12852 17388 12862 17444
rect 13346 17388 13356 17444
rect 13412 17388 13804 17444
rect 13860 17388 13870 17444
rect 14466 17388 14476 17444
rect 14532 17388 14542 17444
rect 19394 17388 19404 17444
rect 19460 17388 19964 17444
rect 20020 17388 20636 17444
rect 20692 17388 21756 17444
rect 21812 17388 21822 17444
rect 22054 17388 22092 17444
rect 22148 17388 22158 17444
rect 22418 17388 22428 17444
rect 22484 17388 23100 17444
rect 23156 17388 23166 17444
rect 5628 17332 5684 17388
rect 14476 17332 14532 17388
rect 3154 17276 3164 17332
rect 3220 17276 3500 17332
rect 3556 17276 4060 17332
rect 4116 17276 5404 17332
rect 5460 17276 5470 17332
rect 5628 17276 7028 17332
rect 7970 17276 7980 17332
rect 8036 17276 14140 17332
rect 14196 17276 14532 17332
rect 15092 17276 15260 17332
rect 15316 17276 19292 17332
rect 19348 17276 19358 17332
rect 21522 17276 21532 17332
rect 21588 17276 21756 17332
rect 21812 17276 21822 17332
rect 6972 17220 7028 17276
rect 15092 17220 15148 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 4386 17164 4396 17220
rect 4452 17164 6804 17220
rect 6934 17164 6972 17220
rect 7028 17164 7038 17220
rect 8418 17164 8428 17220
rect 8484 17164 8522 17220
rect 8866 17164 8876 17220
rect 8932 17164 11564 17220
rect 11620 17164 12684 17220
rect 12740 17164 12750 17220
rect 13990 17164 14028 17220
rect 14084 17164 14094 17220
rect 14466 17164 14476 17220
rect 14532 17164 15148 17220
rect 15922 17164 15932 17220
rect 15988 17164 18396 17220
rect 18452 17164 18508 17220
rect 18564 17164 18574 17220
rect 20850 17164 20860 17220
rect 20916 17164 23548 17220
rect 23604 17164 23660 17220
rect 23716 17164 23726 17220
rect 6748 17108 6804 17164
rect 2006 17052 2044 17108
rect 2100 17052 2110 17108
rect 2594 17052 2604 17108
rect 2660 17052 3164 17108
rect 3220 17052 3230 17108
rect 3332 17052 4956 17108
rect 5012 17052 5022 17108
rect 6738 17052 6748 17108
rect 6804 17052 8540 17108
rect 8596 17052 8606 17108
rect 9090 17052 9100 17108
rect 9156 17052 11956 17108
rect 13570 17052 13580 17108
rect 13636 17052 14252 17108
rect 14308 17052 14588 17108
rect 14644 17052 14654 17108
rect 16146 17052 16156 17108
rect 16212 17052 16492 17108
rect 16548 17052 16558 17108
rect 18722 17052 18732 17108
rect 18788 17052 22092 17108
rect 22148 17052 22158 17108
rect 22642 17052 22652 17108
rect 22708 17052 24332 17108
rect 24388 17052 24398 17108
rect 1894 16940 1932 16996
rect 1988 16940 1998 16996
rect 2678 16940 2716 16996
rect 2772 16940 2782 16996
rect 2716 16884 2772 16940
rect 1698 16828 1708 16884
rect 1764 16828 2772 16884
rect 3332 16772 3388 17052
rect 11900 16996 11956 17052
rect 3714 16940 3724 16996
rect 3780 16940 5068 16996
rect 5124 16940 5134 16996
rect 6290 16940 6300 16996
rect 6356 16940 6524 16996
rect 6580 16940 6590 16996
rect 8306 16940 8316 16996
rect 8372 16940 8764 16996
rect 8820 16940 10220 16996
rect 10276 16940 10286 16996
rect 11890 16940 11900 16996
rect 11956 16940 13468 16996
rect 13524 16940 13534 16996
rect 14018 16940 14028 16996
rect 14084 16940 15372 16996
rect 15428 16940 15438 16996
rect 16034 16940 16044 16996
rect 16100 16940 16660 16996
rect 16930 16940 16940 16996
rect 16996 16940 17388 16996
rect 17444 16940 17724 16996
rect 17780 16940 17790 16996
rect 18498 16940 18508 16996
rect 18564 16940 19068 16996
rect 19124 16940 23996 16996
rect 24052 16940 24780 16996
rect 24836 16940 24846 16996
rect 16604 16884 16660 16940
rect 3826 16828 3836 16884
rect 3892 16828 5964 16884
rect 6020 16828 6030 16884
rect 7522 16828 7532 16884
rect 7588 16828 8204 16884
rect 8260 16828 8270 16884
rect 10546 16828 10556 16884
rect 10612 16828 11228 16884
rect 11284 16828 11294 16884
rect 11778 16828 11788 16884
rect 11844 16828 13692 16884
rect 13748 16828 13758 16884
rect 14690 16828 14700 16884
rect 14756 16828 15596 16884
rect 15652 16828 15662 16884
rect 16230 16828 16268 16884
rect 16324 16828 16334 16884
rect 16566 16828 16604 16884
rect 16660 16828 16670 16884
rect 21634 16828 21644 16884
rect 21700 16828 24388 16884
rect 25218 16828 25228 16884
rect 25284 16828 26460 16884
rect 26516 16828 26526 16884
rect 1026 16716 1036 16772
rect 1092 16716 3388 16772
rect 3714 16716 3724 16772
rect 3780 16716 6412 16772
rect 6468 16716 6478 16772
rect 8614 16716 8652 16772
rect 8708 16716 8718 16772
rect 10882 16716 10892 16772
rect 10948 16716 12124 16772
rect 12180 16716 12190 16772
rect 12786 16716 12796 16772
rect 12852 16716 12964 16772
rect 15222 16716 15260 16772
rect 15316 16716 15326 16772
rect 20514 16716 20524 16772
rect 20580 16716 22652 16772
rect 22708 16716 22718 16772
rect 2258 16604 2268 16660
rect 2324 16604 7868 16660
rect 7924 16604 7934 16660
rect 8082 16604 8092 16660
rect 8148 16604 9660 16660
rect 9716 16604 11340 16660
rect 11396 16604 11406 16660
rect 12226 16604 12236 16660
rect 12292 16604 12572 16660
rect 12628 16604 12638 16660
rect 12908 16548 12964 16716
rect 14242 16604 14252 16660
rect 14308 16604 14812 16660
rect 14868 16604 14878 16660
rect 24332 16548 24388 16828
rect 27458 16716 27468 16772
rect 27524 16716 29484 16772
rect 29540 16716 29550 16772
rect 6850 16492 6860 16548
rect 6916 16492 12684 16548
rect 12740 16492 12750 16548
rect 12908 16492 14140 16548
rect 14196 16492 14476 16548
rect 14532 16492 14542 16548
rect 24332 16492 27468 16548
rect 27524 16492 27534 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 4834 16380 4844 16436
rect 4900 16380 5068 16436
rect 5124 16380 5134 16436
rect 8642 16380 8652 16436
rect 8708 16380 9436 16436
rect 9492 16380 9502 16436
rect 3938 16268 3948 16324
rect 4004 16268 4732 16324
rect 4788 16268 5740 16324
rect 5796 16268 5806 16324
rect 6066 16268 6076 16324
rect 6132 16268 7756 16324
rect 7812 16268 7822 16324
rect 8978 16268 8988 16324
rect 9044 16268 9324 16324
rect 9380 16268 9390 16324
rect 12786 16268 12796 16324
rect 12852 16268 13804 16324
rect 13860 16268 14924 16324
rect 14980 16268 14990 16324
rect 18834 16268 18844 16324
rect 18900 16268 21420 16324
rect 21476 16268 21868 16324
rect 21924 16268 21934 16324
rect 6076 16212 6132 16268
rect 3490 16156 3500 16212
rect 3556 16156 6132 16212
rect 6962 16156 6972 16212
rect 7028 16156 8988 16212
rect 9044 16156 9548 16212
rect 9604 16156 9614 16212
rect 12114 16156 12124 16212
rect 12180 16156 14644 16212
rect 19506 16156 19516 16212
rect 19572 16156 20636 16212
rect 20692 16156 20702 16212
rect 20850 16156 20860 16212
rect 20916 16156 21644 16212
rect 21700 16156 22764 16212
rect 22820 16156 23212 16212
rect 23268 16156 23278 16212
rect 29922 16156 29932 16212
rect 29988 16156 34300 16212
rect 34356 16156 34366 16212
rect 14588 16100 14644 16156
rect 1810 16044 1820 16100
rect 1876 16044 6860 16100
rect 6916 16044 7308 16100
rect 7364 16044 7374 16100
rect 11900 16044 13692 16100
rect 13748 16044 13758 16100
rect 14588 16044 14812 16100
rect 14868 16044 14878 16100
rect 15810 16044 15820 16100
rect 15876 16044 17948 16100
rect 18004 16044 18014 16100
rect 19404 16044 20412 16100
rect 20468 16044 20478 16100
rect 11900 15988 11956 16044
rect 14588 15988 14644 16044
rect 19404 15988 19460 16044
rect 3388 15932 5068 15988
rect 5124 15932 5516 15988
rect 5572 15932 6748 15988
rect 6804 15932 6814 15988
rect 11442 15932 11452 15988
rect 11508 15932 11900 15988
rect 11956 15932 11966 15988
rect 12786 15932 12796 15988
rect 12852 15932 13468 15988
rect 13524 15932 13534 15988
rect 13794 15932 13804 15988
rect 13860 15932 14028 15988
rect 14084 15932 14094 15988
rect 14578 15932 14588 15988
rect 14644 15932 14654 15988
rect 14914 15932 14924 15988
rect 14980 15932 15372 15988
rect 15428 15932 15438 15988
rect 15698 15932 15708 15988
rect 15764 15932 17164 15988
rect 17220 15932 17230 15988
rect 18620 15932 18732 15988
rect 18788 15932 18798 15988
rect 19058 15932 19068 15988
rect 19124 15932 19404 15988
rect 19460 15932 19470 15988
rect 20066 15932 20076 15988
rect 20132 15932 21364 15988
rect 3388 15876 3444 15932
rect 3836 15876 3892 15932
rect 15708 15876 15764 15932
rect 2230 15820 2268 15876
rect 2324 15820 2828 15876
rect 2884 15820 2894 15876
rect 3126 15820 3164 15876
rect 3220 15820 3230 15876
rect 3378 15820 3388 15876
rect 3444 15820 3454 15876
rect 3826 15820 3836 15876
rect 3892 15820 3902 15876
rect 4050 15820 4060 15876
rect 4116 15820 4620 15876
rect 4676 15820 4956 15876
rect 5012 15820 5022 15876
rect 5170 15820 5180 15876
rect 5236 15820 7084 15876
rect 7140 15820 7756 15876
rect 7812 15820 7822 15876
rect 12002 15820 12012 15876
rect 12068 15820 13916 15876
rect 13972 15820 15764 15876
rect 18246 15820 18284 15876
rect 18340 15820 18350 15876
rect 2370 15708 2380 15764
rect 2436 15708 3612 15764
rect 3668 15708 3678 15764
rect 4050 15708 4060 15764
rect 4116 15708 4508 15764
rect 4564 15708 4574 15764
rect 10322 15708 10332 15764
rect 10388 15708 11116 15764
rect 11172 15708 12684 15764
rect 12740 15708 12908 15764
rect 12964 15708 12974 15764
rect 14802 15708 14812 15764
rect 14868 15708 15148 15764
rect 15204 15708 15708 15764
rect 15764 15708 15774 15764
rect 16370 15708 16380 15764
rect 16436 15708 16446 15764
rect 16380 15652 16436 15708
rect 18620 15652 18676 15932
rect 21308 15876 21364 15932
rect 18834 15820 18844 15876
rect 18900 15820 19516 15876
rect 19572 15820 19582 15876
rect 19730 15820 19740 15876
rect 19796 15820 20748 15876
rect 20804 15820 20814 15876
rect 21298 15820 21308 15876
rect 21364 15820 21374 15876
rect 23202 15820 23212 15876
rect 23268 15820 25228 15876
rect 25284 15820 27132 15876
rect 27188 15820 27198 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 7298 15596 7308 15652
rect 7364 15596 12572 15652
rect 12628 15596 14420 15652
rect 14578 15596 14588 15652
rect 14644 15596 17164 15652
rect 17220 15596 17230 15652
rect 18620 15596 19012 15652
rect 20626 15596 20636 15652
rect 20692 15596 21532 15652
rect 21588 15596 21598 15652
rect 14364 15540 14420 15596
rect 3042 15484 3052 15540
rect 3108 15484 3388 15540
rect 5394 15484 5404 15540
rect 5460 15484 7420 15540
rect 7476 15484 7486 15540
rect 8754 15484 8764 15540
rect 8820 15484 9324 15540
rect 9380 15484 9390 15540
rect 9538 15484 9548 15540
rect 9604 15484 9996 15540
rect 10052 15484 10556 15540
rect 10612 15484 10622 15540
rect 11890 15484 11900 15540
rect 11956 15484 13356 15540
rect 13412 15484 13422 15540
rect 14364 15484 14700 15540
rect 14756 15484 14766 15540
rect 16482 15484 16492 15540
rect 16548 15484 16828 15540
rect 16884 15484 17836 15540
rect 17892 15484 17902 15540
rect 3332 15428 3388 15484
rect 18956 15428 19012 15596
rect 19142 15484 19180 15540
rect 19236 15484 19246 15540
rect 19590 15484 19628 15540
rect 19684 15484 19694 15540
rect 20850 15484 20860 15540
rect 20916 15484 22092 15540
rect 22148 15484 22158 15540
rect 24546 15484 24556 15540
rect 24612 15484 24892 15540
rect 24948 15484 28700 15540
rect 28756 15484 30716 15540
rect 30772 15484 30782 15540
rect 3332 15372 3836 15428
rect 3892 15372 3902 15428
rect 4162 15372 4172 15428
rect 4228 15372 5852 15428
rect 5908 15372 5918 15428
rect 6290 15372 6300 15428
rect 6356 15372 12124 15428
rect 12180 15372 12190 15428
rect 13010 15372 13020 15428
rect 13076 15372 15148 15428
rect 17266 15372 17276 15428
rect 17332 15372 18396 15428
rect 18452 15372 18788 15428
rect 18946 15372 18956 15428
rect 19012 15372 19022 15428
rect 22194 15372 22204 15428
rect 22260 15372 22764 15428
rect 22820 15372 22830 15428
rect 23874 15372 23884 15428
rect 23940 15372 24444 15428
rect 24500 15372 24510 15428
rect 24658 15372 24668 15428
rect 24724 15372 25676 15428
rect 25732 15372 26124 15428
rect 26180 15372 26190 15428
rect 28242 15372 28252 15428
rect 28308 15372 30044 15428
rect 30100 15372 31164 15428
rect 31220 15372 36540 15428
rect 36596 15372 36606 15428
rect 15092 15316 15148 15372
rect 18732 15316 18788 15372
rect 1922 15260 1932 15316
rect 1988 15260 4060 15316
rect 4116 15260 4126 15316
rect 4610 15260 4620 15316
rect 4676 15260 6524 15316
rect 6580 15260 6590 15316
rect 8194 15260 8204 15316
rect 8260 15260 8988 15316
rect 9044 15260 10444 15316
rect 10500 15260 10892 15316
rect 10948 15260 10958 15316
rect 11106 15260 11116 15316
rect 11172 15260 11564 15316
rect 11620 15260 12684 15316
rect 12740 15260 12750 15316
rect 13682 15260 13692 15316
rect 13748 15260 14588 15316
rect 14644 15260 14654 15316
rect 15092 15260 15260 15316
rect 15316 15260 17948 15316
rect 18004 15260 18014 15316
rect 18722 15260 18732 15316
rect 18788 15260 18798 15316
rect 18956 15260 20412 15316
rect 20468 15260 20748 15316
rect 20804 15260 20814 15316
rect 21074 15260 21084 15316
rect 21140 15260 21868 15316
rect 21924 15260 21934 15316
rect 22502 15260 22540 15316
rect 22596 15260 22606 15316
rect 23202 15260 23212 15316
rect 23268 15260 23324 15316
rect 23380 15260 23390 15316
rect 25218 15260 25228 15316
rect 25284 15260 26684 15316
rect 26740 15260 26750 15316
rect 27234 15260 27244 15316
rect 27300 15260 28028 15316
rect 28084 15260 29820 15316
rect 29876 15260 31948 15316
rect 32004 15260 32014 15316
rect 3938 15148 3948 15204
rect 4004 15148 7084 15204
rect 7140 15148 7150 15204
rect 7522 15148 7532 15204
rect 7588 15148 8540 15204
rect 8596 15148 8606 15204
rect 10322 15148 10332 15204
rect 10388 15148 12460 15204
rect 12516 15148 12526 15204
rect 13468 15148 15820 15204
rect 15876 15148 15886 15204
rect 16146 15148 16156 15204
rect 16212 15148 16222 15204
rect 13468 15092 13524 15148
rect 16156 15092 16212 15148
rect 18956 15092 19012 15260
rect 19170 15148 19180 15204
rect 19236 15148 19516 15204
rect 19572 15148 20580 15204
rect 25778 15148 25788 15204
rect 25844 15148 26908 15204
rect 26964 15148 27244 15204
rect 27300 15148 27310 15204
rect 28914 15148 28924 15204
rect 28980 15148 30380 15204
rect 30436 15148 32620 15204
rect 32676 15148 33740 15204
rect 33796 15148 33806 15204
rect 20524 15092 20580 15148
rect 4834 15036 4844 15092
rect 4900 15036 7644 15092
rect 7700 15036 11788 15092
rect 11844 15036 11854 15092
rect 13458 15036 13468 15092
rect 13524 15036 13534 15092
rect 15092 15036 16212 15092
rect 18172 15036 19012 15092
rect 20514 15036 20524 15092
rect 20580 15036 20590 15092
rect 26002 15036 26012 15092
rect 26068 15036 26078 15092
rect 15092 14980 15148 15036
rect 5058 14924 5068 14980
rect 5124 14924 6076 14980
rect 6132 14924 6142 14980
rect 8754 14924 8764 14980
rect 8820 14924 9996 14980
rect 10052 14924 10780 14980
rect 10836 14924 10846 14980
rect 14140 14924 14476 14980
rect 14532 14924 15148 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 14140 14868 14196 14924
rect 3378 14812 3388 14868
rect 3444 14812 4284 14868
rect 4340 14812 4350 14868
rect 5180 14812 14196 14868
rect 5180 14756 5236 14812
rect 3826 14700 3836 14756
rect 3892 14700 5236 14756
rect 5394 14700 5404 14756
rect 5460 14700 5740 14756
rect 5796 14700 5806 14756
rect 7942 14700 7980 14756
rect 8036 14700 8046 14756
rect 9314 14700 9324 14756
rect 9380 14700 9772 14756
rect 9828 14700 9838 14756
rect 11638 14700 11676 14756
rect 11732 14700 11742 14756
rect 14998 14700 15036 14756
rect 15092 14700 15102 14756
rect 1922 14588 1932 14644
rect 1988 14588 2156 14644
rect 2212 14588 3388 14644
rect 5506 14588 5516 14644
rect 5572 14588 13468 14644
rect 13524 14588 13534 14644
rect 14130 14588 14140 14644
rect 14196 14588 14812 14644
rect 14868 14588 14878 14644
rect 15894 14588 15932 14644
rect 15988 14588 15998 14644
rect 3332 14532 3388 14588
rect 3332 14476 7980 14532
rect 8036 14476 8046 14532
rect 14018 14476 14028 14532
rect 14084 14476 15036 14532
rect 15092 14476 16268 14532
rect 16324 14476 16334 14532
rect 18172 14420 18228 15036
rect 18386 14924 18396 14980
rect 18452 14924 18620 14980
rect 18676 14924 18686 14980
rect 21746 14924 21756 14980
rect 21812 14924 22764 14980
rect 22820 14924 22830 14980
rect 23762 14924 23772 14980
rect 23828 14924 25452 14980
rect 25508 14924 25518 14980
rect 26012 14868 26068 15036
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 22866 14812 22876 14868
rect 22932 14812 23996 14868
rect 24052 14812 24062 14868
rect 25330 14812 25340 14868
rect 25396 14812 26068 14868
rect 19394 14700 19404 14756
rect 19460 14700 20188 14756
rect 20244 14700 20254 14756
rect 22978 14700 22988 14756
rect 23044 14700 23772 14756
rect 23828 14700 23838 14756
rect 21942 14588 21980 14644
rect 22036 14588 22046 14644
rect 27458 14588 27468 14644
rect 27524 14588 28028 14644
rect 28084 14588 42140 14644
rect 42196 14588 42206 14644
rect 19506 14476 19516 14532
rect 19572 14476 20076 14532
rect 20132 14476 20142 14532
rect 20402 14476 20412 14532
rect 20468 14476 20636 14532
rect 20692 14476 20702 14532
rect 26852 14476 32844 14532
rect 32900 14476 32910 14532
rect 26852 14420 26908 14476
rect 3490 14364 3500 14420
rect 3556 14364 7420 14420
rect 7476 14364 7486 14420
rect 12562 14364 12572 14420
rect 12628 14364 13356 14420
rect 13412 14364 13422 14420
rect 14578 14364 14588 14420
rect 14644 14364 18228 14420
rect 19180 14364 19292 14420
rect 19348 14364 21980 14420
rect 22036 14364 22046 14420
rect 26002 14364 26012 14420
rect 26068 14364 26908 14420
rect 29932 14364 33292 14420
rect 33348 14364 33358 14420
rect 19180 14308 19236 14364
rect 29932 14308 29988 14364
rect 3574 14252 3612 14308
rect 3668 14252 3678 14308
rect 4050 14252 4060 14308
rect 4116 14252 4284 14308
rect 4340 14252 4396 14308
rect 4452 14252 4462 14308
rect 4946 14252 4956 14308
rect 5012 14252 5852 14308
rect 5908 14252 6076 14308
rect 6132 14252 6142 14308
rect 6402 14252 6412 14308
rect 6468 14252 6692 14308
rect 6962 14252 6972 14308
rect 7028 14252 7196 14308
rect 7252 14252 7262 14308
rect 8082 14252 8092 14308
rect 8148 14252 8652 14308
rect 8708 14252 9660 14308
rect 9716 14252 9726 14308
rect 11218 14252 11228 14308
rect 11284 14252 11788 14308
rect 11844 14252 15148 14308
rect 17266 14252 17276 14308
rect 17332 14252 17836 14308
rect 17892 14252 17902 14308
rect 18162 14252 18172 14308
rect 18228 14252 19236 14308
rect 19394 14252 19404 14308
rect 19460 14252 20300 14308
rect 20356 14252 20366 14308
rect 20626 14252 20636 14308
rect 20692 14252 22204 14308
rect 22260 14252 22270 14308
rect 26674 14252 26684 14308
rect 26740 14252 27132 14308
rect 27188 14252 27198 14308
rect 27542 14252 27580 14308
rect 27636 14252 27646 14308
rect 28802 14252 28812 14308
rect 28868 14252 29484 14308
rect 29540 14252 29932 14308
rect 29988 14252 29998 14308
rect 30930 14252 30940 14308
rect 30996 14252 31612 14308
rect 31668 14252 32396 14308
rect 32452 14252 32462 14308
rect 6636 14196 6692 14252
rect 15092 14196 15148 14252
rect 2258 14140 2268 14196
rect 2324 14140 3836 14196
rect 3892 14140 4284 14196
rect 4340 14140 4350 14196
rect 6626 14140 6636 14196
rect 6692 14140 6702 14196
rect 11676 14140 13244 14196
rect 13300 14140 13580 14196
rect 13636 14140 13646 14196
rect 15092 14140 15260 14196
rect 15316 14140 16716 14196
rect 16772 14140 16782 14196
rect 17042 14140 17052 14196
rect 17108 14140 18060 14196
rect 18116 14140 18508 14196
rect 18564 14140 18574 14196
rect 11676 14084 11732 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 6738 14028 6748 14084
rect 6804 14028 7868 14084
rect 7924 14028 11116 14084
rect 11172 14028 11732 14084
rect 12002 14028 12012 14084
rect 12068 14028 16380 14084
rect 16436 14028 16446 14084
rect 19058 14028 19068 14084
rect 19124 14028 19516 14084
rect 19572 14028 19582 14084
rect 20402 14028 20412 14084
rect 20468 14028 21756 14084
rect 21812 14028 21980 14084
rect 22036 14028 23100 14084
rect 23156 14028 23166 14084
rect 4946 13916 4956 13972
rect 5012 13916 5022 13972
rect 8540 13916 8876 13972
rect 8932 13916 8942 13972
rect 9874 13916 9884 13972
rect 9940 13916 9996 13972
rect 10052 13916 10062 13972
rect 10210 13916 10220 13972
rect 10276 13916 10892 13972
rect 10948 13916 10958 13972
rect 12450 13916 12460 13972
rect 12516 13916 15148 13972
rect 15204 13916 16604 13972
rect 16660 13916 16670 13972
rect 18722 13916 18732 13972
rect 18788 13916 21420 13972
rect 21476 13916 21486 13972
rect 22082 13916 22092 13972
rect 22148 13916 23324 13972
rect 23380 13916 24556 13972
rect 24612 13916 24622 13972
rect 26338 13916 26348 13972
rect 26404 13916 28140 13972
rect 28196 13916 28206 13972
rect 29026 13916 29036 13972
rect 29092 13916 31948 13972
rect 32004 13916 32172 13972
rect 32228 13916 34748 13972
rect 34804 13916 34814 13972
rect 4956 13860 5012 13916
rect 8540 13860 8596 13916
rect 4956 13804 7308 13860
rect 7364 13804 7374 13860
rect 8194 13804 8204 13860
rect 8260 13804 8596 13860
rect 8754 13804 8764 13860
rect 8820 13804 10108 13860
rect 10164 13804 10174 13860
rect 12786 13804 12796 13860
rect 12852 13804 15820 13860
rect 15876 13804 15886 13860
rect 18834 13804 18844 13860
rect 18900 13804 20524 13860
rect 20580 13804 20590 13860
rect 22642 13804 22652 13860
rect 22708 13804 22718 13860
rect 23874 13804 23884 13860
rect 23940 13804 24444 13860
rect 24500 13804 24510 13860
rect 25554 13804 25564 13860
rect 25620 13804 26572 13860
rect 26628 13804 26638 13860
rect 31714 13804 31724 13860
rect 31780 13804 32284 13860
rect 32340 13804 32350 13860
rect 22652 13748 22708 13804
rect 4834 13692 4844 13748
rect 4900 13692 5180 13748
rect 5236 13692 5246 13748
rect 5590 13692 5628 13748
rect 5684 13692 5694 13748
rect 7858 13692 7868 13748
rect 7924 13692 13356 13748
rect 13412 13692 13422 13748
rect 13570 13692 13580 13748
rect 13636 13692 15596 13748
rect 15652 13692 15662 13748
rect 16706 13692 16716 13748
rect 16772 13692 18620 13748
rect 18676 13692 18686 13748
rect 19170 13692 19180 13748
rect 19236 13692 22708 13748
rect 26002 13692 26012 13748
rect 26068 13692 27132 13748
rect 27188 13692 27198 13748
rect 28802 13692 28812 13748
rect 28868 13692 29820 13748
rect 29876 13692 29886 13748
rect 1922 13580 1932 13636
rect 1988 13580 3164 13636
rect 3220 13580 3230 13636
rect 4050 13580 4060 13636
rect 4116 13580 7308 13636
rect 7364 13580 7374 13636
rect 14914 13580 14924 13636
rect 14980 13580 17892 13636
rect 18162 13580 18172 13636
rect 18228 13580 19068 13636
rect 19124 13580 22652 13636
rect 22708 13580 22718 13636
rect 26786 13580 26796 13636
rect 26852 13580 29372 13636
rect 29428 13580 31164 13636
rect 31220 13580 32620 13636
rect 32676 13580 33404 13636
rect 33460 13580 33470 13636
rect 2034 13468 2044 13524
rect 2100 13468 3724 13524
rect 3780 13468 4844 13524
rect 4900 13468 4910 13524
rect 6402 13468 6412 13524
rect 6468 13468 10556 13524
rect 10612 13468 10622 13524
rect 11554 13468 11564 13524
rect 11620 13468 12460 13524
rect 12516 13468 12526 13524
rect 12674 13468 12684 13524
rect 12740 13468 14476 13524
rect 14532 13468 14542 13524
rect 14802 13468 14812 13524
rect 14868 13468 15372 13524
rect 15428 13468 15820 13524
rect 15876 13468 15886 13524
rect 17836 13412 17892 13580
rect 18050 13468 18060 13524
rect 18116 13468 19628 13524
rect 19684 13468 19694 13524
rect 22194 13468 22204 13524
rect 22260 13468 22764 13524
rect 22820 13468 22830 13524
rect 23314 13468 23324 13524
rect 23380 13468 24556 13524
rect 24612 13468 26348 13524
rect 26404 13468 26414 13524
rect 26674 13468 26684 13524
rect 26740 13468 27020 13524
rect 27076 13468 27468 13524
rect 27524 13468 27534 13524
rect 9874 13356 9884 13412
rect 9940 13356 10220 13412
rect 10276 13356 10286 13412
rect 12786 13356 12796 13412
rect 12852 13356 15260 13412
rect 15316 13356 15326 13412
rect 17836 13356 19292 13412
rect 19348 13356 19358 13412
rect 19618 13356 19628 13412
rect 19684 13356 19852 13412
rect 19908 13356 19918 13412
rect 22642 13356 22652 13412
rect 22708 13356 24332 13412
rect 24388 13356 24398 13412
rect 24658 13356 24668 13412
rect 24724 13356 25564 13412
rect 25620 13356 25630 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 3826 13244 3836 13300
rect 3892 13244 4060 13300
rect 4116 13244 4126 13300
rect 14914 13244 14924 13300
rect 14980 13244 15036 13300
rect 15092 13244 15102 13300
rect 19506 13244 19516 13300
rect 19572 13244 20860 13300
rect 20916 13244 20926 13300
rect 21074 13244 21084 13300
rect 21140 13244 22876 13300
rect 22932 13244 23548 13300
rect 23604 13244 28140 13300
rect 28196 13244 28476 13300
rect 28532 13244 28542 13300
rect 3042 13132 3052 13188
rect 3108 13132 6860 13188
rect 6916 13132 6926 13188
rect 9090 13132 9100 13188
rect 9156 13132 11676 13188
rect 11732 13132 14364 13188
rect 14420 13132 14430 13188
rect 16818 13132 16828 13188
rect 16884 13132 17388 13188
rect 17444 13132 17454 13188
rect 17938 13132 17948 13188
rect 18004 13132 22540 13188
rect 22596 13132 25564 13188
rect 25620 13132 25630 13188
rect 32162 13132 32172 13188
rect 32228 13132 32396 13188
rect 32452 13132 32462 13188
rect 3714 13020 3724 13076
rect 3780 13020 6972 13076
rect 7028 13020 7038 13076
rect 7186 13020 7196 13076
rect 7252 13020 8204 13076
rect 8260 13020 8270 13076
rect 14578 13020 14588 13076
rect 14644 13020 24220 13076
rect 24276 13020 24286 13076
rect 24434 13020 24444 13076
rect 24500 13020 27244 13076
rect 27300 13020 27310 13076
rect 5964 12964 6020 13020
rect 6972 12964 7028 13020
rect 2930 12908 2940 12964
rect 2996 12908 3388 12964
rect 3444 12908 4676 12964
rect 4834 12908 4844 12964
rect 4900 12908 5068 12964
rect 5124 12908 5134 12964
rect 5366 12908 5404 12964
rect 5460 12908 5470 12964
rect 5954 12908 5964 12964
rect 6020 12908 6030 12964
rect 6972 12908 8428 12964
rect 8484 12908 8494 12964
rect 13346 12908 13356 12964
rect 13412 12908 14812 12964
rect 14868 12908 14878 12964
rect 20066 12908 20076 12964
rect 20132 12908 21196 12964
rect 21252 12908 21262 12964
rect 22754 12908 22764 12964
rect 22820 12908 22830 12964
rect 23090 12908 23100 12964
rect 23156 12908 23166 12964
rect 4620 12852 4676 12908
rect 22764 12852 22820 12908
rect 23100 12852 23156 12908
rect 2258 12796 2268 12852
rect 2324 12796 2492 12852
rect 2548 12796 2558 12852
rect 3266 12796 3276 12852
rect 3332 12796 4396 12852
rect 4452 12796 4462 12852
rect 4620 12796 6972 12852
rect 7028 12796 8372 12852
rect 8530 12796 8540 12852
rect 8596 12796 8876 12852
rect 8932 12796 13692 12852
rect 13748 12796 19740 12852
rect 19796 12796 22540 12852
rect 22596 12796 22820 12852
rect 22876 12796 23156 12852
rect 24220 12852 24276 13020
rect 26450 12908 26460 12964
rect 26516 12908 27916 12964
rect 27972 12908 27982 12964
rect 24220 12796 27468 12852
rect 27524 12796 27692 12852
rect 27748 12796 27758 12852
rect 30258 12796 30268 12852
rect 30324 12796 31276 12852
rect 31332 12796 31342 12852
rect 35522 12796 35532 12852
rect 35588 12796 36932 12852
rect 8316 12740 8372 12796
rect 3938 12684 3948 12740
rect 4004 12684 6748 12740
rect 6804 12684 6814 12740
rect 7410 12684 7420 12740
rect 7476 12684 8092 12740
rect 8148 12684 8158 12740
rect 8316 12684 10220 12740
rect 10276 12684 10286 12740
rect 10882 12684 10892 12740
rect 10948 12684 22316 12740
rect 22372 12684 22382 12740
rect 22876 12628 22932 12796
rect 36876 12740 36932 12796
rect 23024 12684 23100 12740
rect 23156 12684 24556 12740
rect 24612 12684 24622 12740
rect 24780 12684 30716 12740
rect 30772 12684 30782 12740
rect 34290 12684 34300 12740
rect 34356 12684 35084 12740
rect 35140 12684 36428 12740
rect 36484 12684 36652 12740
rect 36708 12684 36718 12740
rect 36876 12684 40572 12740
rect 40628 12684 40638 12740
rect 24780 12628 24836 12684
rect 30268 12628 30324 12684
rect 3714 12572 3724 12628
rect 3780 12572 5068 12628
rect 5124 12572 6412 12628
rect 6468 12572 6478 12628
rect 7522 12572 7532 12628
rect 7588 12572 8988 12628
rect 9044 12572 9054 12628
rect 15586 12572 15596 12628
rect 15652 12572 16268 12628
rect 16324 12572 16940 12628
rect 16996 12572 17006 12628
rect 21970 12572 21980 12628
rect 22036 12572 24836 12628
rect 25666 12572 25676 12628
rect 25732 12572 26908 12628
rect 26964 12572 28868 12628
rect 30258 12572 30268 12628
rect 30324 12572 30334 12628
rect 33618 12572 33628 12628
rect 33684 12572 34748 12628
rect 34804 12572 34814 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 28812 12516 28868 12572
rect 1922 12460 1932 12516
rect 1988 12460 7196 12516
rect 7252 12460 7262 12516
rect 15810 12460 15820 12516
rect 15876 12460 18284 12516
rect 18340 12460 18350 12516
rect 19058 12460 19068 12516
rect 19124 12460 19180 12516
rect 19236 12460 19246 12516
rect 22082 12460 22092 12516
rect 22148 12460 22540 12516
rect 22596 12460 22606 12516
rect 23212 12460 23772 12516
rect 23828 12460 23996 12516
rect 24052 12460 24062 12516
rect 26338 12460 26348 12516
rect 26404 12460 26414 12516
rect 26786 12460 26796 12516
rect 26852 12460 28364 12516
rect 28420 12460 28430 12516
rect 28802 12460 28812 12516
rect 28868 12460 32956 12516
rect 33012 12460 33022 12516
rect 34178 12460 34188 12516
rect 34244 12460 34972 12516
rect 35028 12460 35038 12516
rect 35858 12460 35868 12516
rect 35924 12460 42028 12516
rect 42084 12460 42812 12516
rect 42868 12460 42878 12516
rect 23212 12404 23268 12460
rect 2594 12348 2604 12404
rect 2660 12348 3836 12404
rect 3892 12348 3902 12404
rect 4050 12348 4060 12404
rect 4116 12348 5180 12404
rect 5236 12348 7084 12404
rect 7140 12348 7150 12404
rect 7494 12348 7532 12404
rect 7588 12348 7598 12404
rect 9090 12348 9100 12404
rect 9156 12348 14588 12404
rect 14644 12348 14654 12404
rect 16370 12348 16380 12404
rect 16436 12348 16940 12404
rect 16996 12348 17006 12404
rect 23202 12348 23212 12404
rect 23268 12348 23278 12404
rect 2146 12236 2156 12292
rect 2212 12236 3948 12292
rect 4004 12236 4014 12292
rect 4162 12236 4172 12292
rect 4228 12236 4732 12292
rect 4788 12236 4844 12292
rect 4900 12236 7756 12292
rect 7812 12236 7822 12292
rect 10994 12236 11004 12292
rect 11060 12236 11564 12292
rect 11620 12236 11630 12292
rect 15922 12236 15932 12292
rect 15988 12236 16268 12292
rect 16324 12236 16334 12292
rect 20514 12236 20524 12292
rect 20580 12236 20860 12292
rect 20916 12236 21644 12292
rect 21700 12236 22316 12292
rect 22372 12236 22382 12292
rect 2604 12180 2660 12236
rect 23436 12180 23492 12404
rect 23548 12348 23558 12404
rect 24994 12348 25004 12404
rect 25060 12348 25788 12404
rect 25844 12348 25854 12404
rect 26348 12292 26404 12460
rect 23622 12236 23660 12292
rect 23716 12236 23726 12292
rect 26348 12236 27468 12292
rect 27524 12236 27534 12292
rect 28802 12236 28812 12292
rect 28868 12236 32172 12292
rect 32228 12236 32732 12292
rect 32788 12236 33964 12292
rect 34020 12236 35084 12292
rect 35140 12236 35150 12292
rect 2594 12124 2604 12180
rect 2660 12124 2670 12180
rect 2818 12124 2828 12180
rect 2884 12124 3164 12180
rect 3220 12124 3724 12180
rect 3780 12124 3790 12180
rect 18162 12124 18172 12180
rect 18228 12124 19628 12180
rect 19684 12124 22988 12180
rect 23044 12124 23054 12180
rect 23426 12124 23436 12180
rect 23492 12124 23502 12180
rect 24070 12124 24108 12180
rect 24164 12124 24174 12180
rect 27010 12124 27020 12180
rect 27076 12124 30156 12180
rect 30212 12124 30222 12180
rect 30604 12124 32844 12180
rect 32900 12124 33292 12180
rect 33348 12124 33358 12180
rect 30604 12068 30660 12124
rect 3826 12012 3836 12068
rect 3892 12012 4284 12068
rect 4340 12012 4350 12068
rect 6290 12012 6300 12068
rect 6356 12012 11676 12068
rect 11732 12012 11742 12068
rect 12562 12012 12572 12068
rect 12628 12012 14588 12068
rect 14644 12012 14654 12068
rect 21970 12012 21980 12068
rect 22036 12012 23100 12068
rect 23156 12012 23166 12068
rect 23314 12012 23324 12068
rect 23380 12012 23418 12068
rect 26898 12012 26908 12068
rect 26964 12012 28364 12068
rect 28420 12012 28430 12068
rect 29148 12012 30604 12068
rect 30660 12012 30670 12068
rect 30930 12012 30940 12068
rect 30996 12012 31836 12068
rect 31892 12012 36540 12068
rect 36596 12012 36606 12068
rect 36754 12012 36764 12068
rect 36820 12012 37884 12068
rect 37940 12012 37950 12068
rect 11676 11956 11732 12012
rect 29148 11956 29204 12012
rect 2482 11900 2492 11956
rect 2548 11900 3500 11956
rect 3556 11900 3566 11956
rect 5730 11900 5740 11956
rect 5796 11900 8764 11956
rect 8820 11900 8830 11956
rect 11676 11900 16716 11956
rect 16772 11900 16782 11956
rect 21746 11900 21756 11956
rect 21812 11900 24444 11956
rect 24500 11900 24510 11956
rect 26758 11900 26796 11956
rect 26852 11900 26862 11956
rect 27794 11900 27804 11956
rect 27860 11900 28252 11956
rect 28308 11900 29204 11956
rect 29362 11900 29372 11956
rect 29428 11900 30828 11956
rect 30884 11900 30894 11956
rect 31490 11900 31500 11956
rect 31556 11900 33628 11956
rect 33684 11900 33694 11956
rect 33954 11900 33964 11956
rect 34020 11900 35532 11956
rect 35588 11900 35598 11956
rect 3500 11844 3556 11900
rect 3500 11788 3724 11844
rect 3780 11788 3790 11844
rect 6738 11788 6748 11844
rect 6804 11788 6814 11844
rect 6962 11788 6972 11844
rect 7028 11788 7644 11844
rect 7700 11788 7710 11844
rect 9314 11788 9324 11844
rect 9380 11788 9390 11844
rect 9660 11788 9772 11844
rect 9828 11788 9838 11844
rect 9986 11788 9996 11844
rect 10052 11788 10220 11844
rect 10276 11788 12236 11844
rect 12292 11788 12302 11844
rect 20402 11788 20412 11844
rect 20468 11788 21868 11844
rect 21924 11788 21934 11844
rect 22642 11788 22652 11844
rect 22708 11788 24892 11844
rect 24948 11788 24958 11844
rect 27206 11788 27244 11844
rect 27300 11788 27310 11844
rect 30342 11788 30380 11844
rect 30436 11788 30446 11844
rect 37426 11788 37436 11844
rect 37492 11788 37996 11844
rect 38052 11788 38062 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 6748 11732 6804 11788
rect 9324 11732 9380 11788
rect 9660 11732 9716 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 1810 11676 1820 11732
rect 1876 11676 3276 11732
rect 3332 11676 3342 11732
rect 4834 11676 4844 11732
rect 4900 11676 5852 11732
rect 5908 11676 5918 11732
rect 6748 11676 7196 11732
rect 7252 11676 7262 11732
rect 8306 11676 8316 11732
rect 8372 11676 9716 11732
rect 9874 11676 9884 11732
rect 9940 11676 22708 11732
rect 23538 11676 23548 11732
rect 23604 11676 24556 11732
rect 24612 11676 25676 11732
rect 25732 11676 25742 11732
rect 31714 11676 31724 11732
rect 31780 11676 32396 11732
rect 32452 11676 32462 11732
rect 35746 11676 35756 11732
rect 35812 11676 36204 11732
rect 36260 11676 36988 11732
rect 37044 11676 37772 11732
rect 37828 11676 37838 11732
rect 3388 11564 6188 11620
rect 6244 11564 6254 11620
rect 9314 11564 9324 11620
rect 9380 11564 10668 11620
rect 10724 11564 10734 11620
rect 14914 11564 14924 11620
rect 14980 11564 15036 11620
rect 15092 11564 15102 11620
rect 15362 11564 15372 11620
rect 15428 11564 18060 11620
rect 18116 11564 18620 11620
rect 18676 11564 18686 11620
rect 3388 11508 3444 11564
rect 22652 11508 22708 11676
rect 23426 11564 23436 11620
rect 23492 11564 23660 11620
rect 23716 11564 23726 11620
rect 23874 11564 23884 11620
rect 23940 11564 25116 11620
rect 25172 11564 25788 11620
rect 25844 11564 28700 11620
rect 28756 11564 29596 11620
rect 29652 11564 29662 11620
rect 29810 11564 29820 11620
rect 29876 11564 32060 11620
rect 32116 11564 32126 11620
rect 3378 11452 3388 11508
rect 3444 11452 3454 11508
rect 5740 11452 9212 11508
rect 9268 11452 9772 11508
rect 9828 11452 10220 11508
rect 10276 11452 10286 11508
rect 16818 11452 16828 11508
rect 16884 11452 17500 11508
rect 17556 11452 21812 11508
rect 22652 11452 25340 11508
rect 25396 11452 26684 11508
rect 26740 11452 26750 11508
rect 28578 11452 28588 11508
rect 28644 11452 30884 11508
rect 31042 11452 31052 11508
rect 31108 11452 31500 11508
rect 31556 11452 32620 11508
rect 32676 11452 32686 11508
rect 5740 11396 5796 11452
rect 1138 11340 1148 11396
rect 1204 11340 5068 11396
rect 5124 11340 5516 11396
rect 5572 11340 5582 11396
rect 5730 11340 5740 11396
rect 5796 11340 5834 11396
rect 6598 11340 6636 11396
rect 6692 11340 6702 11396
rect 8866 11340 8876 11396
rect 8932 11340 10108 11396
rect 10164 11340 10174 11396
rect 11218 11340 11228 11396
rect 11284 11340 11452 11396
rect 11508 11340 12460 11396
rect 12516 11340 12526 11396
rect 16258 11340 16268 11396
rect 16324 11340 17388 11396
rect 17444 11340 17454 11396
rect 19394 11340 19404 11396
rect 19460 11340 21532 11396
rect 21588 11340 21598 11396
rect 21756 11284 21812 11452
rect 30828 11396 30884 11452
rect 22194 11340 22204 11396
rect 22260 11340 23436 11396
rect 23492 11340 23996 11396
rect 24052 11340 25004 11396
rect 25060 11340 25070 11396
rect 26002 11340 26012 11396
rect 26068 11340 27356 11396
rect 27412 11340 27422 11396
rect 29810 11340 29820 11396
rect 29876 11340 29932 11396
rect 29988 11340 29998 11396
rect 30828 11340 33180 11396
rect 33236 11340 33628 11396
rect 33684 11340 33694 11396
rect 37650 11340 37660 11396
rect 37716 11340 38668 11396
rect 38724 11340 38734 11396
rect 38994 11340 39004 11396
rect 39060 11340 39676 11396
rect 39732 11340 39742 11396
rect 3154 11228 3164 11284
rect 3220 11228 6524 11284
rect 6580 11228 6590 11284
rect 12562 11228 12572 11284
rect 12628 11228 14700 11284
rect 14756 11228 14766 11284
rect 15698 11228 15708 11284
rect 15764 11228 16156 11284
rect 16212 11228 16222 11284
rect 17490 11228 17500 11284
rect 17556 11228 18788 11284
rect 21756 11228 24892 11284
rect 24948 11228 31052 11284
rect 31108 11228 31118 11284
rect 34626 11228 34636 11284
rect 34692 11228 37548 11284
rect 37604 11228 37614 11284
rect 18732 11172 18788 11228
rect 5170 11116 5180 11172
rect 5236 11116 7532 11172
rect 7588 11116 7598 11172
rect 9734 11116 9772 11172
rect 9828 11116 9838 11172
rect 9986 11116 9996 11172
rect 10052 11116 10108 11172
rect 10164 11116 10174 11172
rect 11666 11116 11676 11172
rect 11732 11116 11742 11172
rect 12450 11116 12460 11172
rect 12516 11116 14028 11172
rect 14084 11116 14094 11172
rect 16482 11116 16492 11172
rect 16548 11116 17276 11172
rect 17332 11116 17612 11172
rect 17668 11116 17836 11172
rect 17892 11116 17902 11172
rect 18722 11116 18732 11172
rect 18788 11116 19852 11172
rect 19908 11116 20524 11172
rect 20580 11116 20590 11172
rect 21410 11116 21420 11172
rect 21476 11116 22764 11172
rect 22820 11116 22830 11172
rect 22988 11116 25228 11172
rect 25284 11116 25294 11172
rect 25890 11116 25900 11172
rect 25956 11116 26124 11172
rect 26180 11116 26572 11172
rect 26628 11116 26638 11172
rect 26786 11116 26796 11172
rect 0 11060 800 11088
rect 11676 11060 11732 11116
rect 22988 11060 23044 11116
rect 0 11004 1820 11060
rect 1876 11004 1932 11060
rect 1988 11004 1998 11060
rect 6626 11004 6636 11060
rect 6692 11004 8204 11060
rect 8260 11004 8270 11060
rect 9314 11004 9324 11060
rect 9380 11004 13692 11060
rect 13748 11004 14252 11060
rect 14308 11004 16212 11060
rect 18610 11004 18620 11060
rect 18676 11004 19628 11060
rect 19684 11004 19694 11060
rect 21186 11004 21196 11060
rect 21252 11004 21868 11060
rect 21924 11004 23044 11060
rect 26852 11060 26908 11172
rect 27346 11116 27356 11172
rect 27412 11116 29820 11172
rect 29876 11116 29886 11172
rect 30370 11116 30380 11172
rect 30436 11116 30716 11172
rect 30772 11116 32060 11172
rect 32116 11116 32126 11172
rect 32834 11116 32844 11172
rect 32900 11116 33516 11172
rect 33572 11116 33582 11172
rect 26852 11004 27300 11060
rect 27458 11004 27468 11060
rect 27524 11004 29484 11060
rect 29540 11004 29550 11060
rect 0 10976 800 11004
rect 4386 10892 4396 10948
rect 4452 10892 6860 10948
rect 6916 10892 6926 10948
rect 15138 10892 15148 10948
rect 15204 10892 15820 10948
rect 15876 10892 15886 10948
rect 16156 10836 16212 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 20188 10892 27188 10948
rect 20188 10836 20244 10892
rect 4498 10780 4508 10836
rect 4564 10780 6076 10836
rect 6132 10780 6142 10836
rect 6514 10780 6524 10836
rect 6580 10780 8428 10836
rect 8484 10780 9100 10836
rect 9156 10780 9996 10836
rect 10052 10780 11004 10836
rect 11060 10780 11070 10836
rect 14802 10780 14812 10836
rect 14868 10780 15372 10836
rect 15428 10780 15438 10836
rect 16146 10780 16156 10836
rect 16212 10780 18508 10836
rect 18564 10780 20244 10836
rect 23874 10780 23884 10836
rect 23940 10780 24108 10836
rect 24164 10780 24174 10836
rect 24556 10780 26908 10836
rect 26964 10780 26974 10836
rect 5618 10668 5628 10724
rect 5684 10668 7308 10724
rect 7364 10668 7374 10724
rect 7644 10668 11340 10724
rect 11396 10668 11406 10724
rect 17042 10668 17052 10724
rect 17108 10668 22092 10724
rect 22148 10668 22158 10724
rect 3602 10556 3612 10612
rect 3668 10556 4172 10612
rect 4228 10556 4238 10612
rect 5730 10556 5740 10612
rect 5796 10556 6188 10612
rect 6244 10556 7420 10612
rect 7476 10556 7486 10612
rect 7644 10500 7700 10668
rect 9762 10556 9772 10612
rect 9828 10556 10332 10612
rect 10388 10556 10398 10612
rect 11218 10556 11228 10612
rect 11284 10556 16380 10612
rect 16436 10556 16446 10612
rect 18470 10556 18508 10612
rect 18564 10556 18574 10612
rect 19170 10556 19180 10612
rect 19236 10556 22204 10612
rect 22260 10556 22270 10612
rect 6738 10444 6748 10500
rect 6804 10444 7532 10500
rect 7588 10444 7700 10500
rect 10780 10444 11564 10500
rect 11620 10444 11630 10500
rect 11890 10444 11900 10500
rect 11956 10444 14924 10500
rect 14980 10444 14990 10500
rect 16594 10444 16604 10500
rect 16660 10444 20524 10500
rect 20580 10444 23100 10500
rect 23156 10444 23166 10500
rect 10780 10388 10836 10444
rect 24556 10388 24612 10780
rect 27132 10724 27188 10892
rect 27244 10836 27300 11004
rect 33394 10892 33404 10948
rect 33460 10892 33628 10948
rect 33684 10892 37660 10948
rect 37716 10892 37726 10948
rect 27244 10780 28588 10836
rect 28644 10780 28654 10836
rect 34514 10780 34524 10836
rect 34580 10780 36092 10836
rect 36148 10780 36158 10836
rect 38210 10780 38220 10836
rect 38276 10780 39228 10836
rect 39284 10780 39294 10836
rect 39554 10780 39564 10836
rect 39620 10780 40236 10836
rect 40292 10780 40572 10836
rect 40628 10780 40638 10836
rect 25218 10668 25228 10724
rect 25284 10668 26236 10724
rect 26292 10668 26796 10724
rect 26852 10668 26862 10724
rect 27132 10668 27468 10724
rect 27524 10668 27534 10724
rect 29250 10668 29260 10724
rect 29316 10668 30268 10724
rect 30324 10668 30334 10724
rect 36866 10668 36876 10724
rect 36932 10668 39116 10724
rect 39172 10668 39182 10724
rect 34178 10556 34188 10612
rect 34244 10556 35532 10612
rect 35588 10556 35598 10612
rect 37986 10556 37996 10612
rect 38052 10556 38556 10612
rect 38612 10556 39004 10612
rect 39060 10556 39070 10612
rect 39778 10556 39788 10612
rect 39844 10556 40124 10612
rect 40180 10556 41356 10612
rect 41412 10556 41422 10612
rect 26786 10444 26796 10500
rect 26852 10444 27356 10500
rect 27412 10444 27422 10500
rect 31826 10444 31836 10500
rect 31892 10444 32396 10500
rect 32452 10444 32462 10500
rect 37762 10444 37772 10500
rect 37828 10444 41804 10500
rect 41860 10444 41870 10500
rect 4050 10332 4060 10388
rect 4116 10332 5292 10388
rect 5348 10332 5358 10388
rect 6178 10332 6188 10388
rect 6244 10332 8316 10388
rect 8372 10332 8382 10388
rect 10210 10332 10220 10388
rect 10276 10332 10780 10388
rect 10836 10332 10846 10388
rect 11330 10332 11340 10388
rect 11396 10332 16268 10388
rect 16324 10332 18060 10388
rect 18116 10332 18126 10388
rect 22754 10332 22764 10388
rect 22820 10332 24556 10388
rect 24612 10332 24622 10388
rect 25778 10332 25788 10388
rect 25844 10332 29708 10388
rect 29764 10332 29774 10388
rect 36082 10332 36092 10388
rect 36148 10332 38556 10388
rect 38612 10332 39676 10388
rect 39732 10332 41972 10388
rect 41916 10276 41972 10332
rect 3602 10220 3612 10276
rect 3668 10220 3948 10276
rect 4004 10220 4014 10276
rect 11330 10220 11340 10276
rect 11396 10220 23548 10276
rect 23604 10220 23614 10276
rect 24994 10220 25004 10276
rect 25060 10220 26684 10276
rect 26740 10220 26750 10276
rect 37436 10220 39228 10276
rect 39284 10220 39788 10276
rect 39844 10220 39854 10276
rect 41906 10220 41916 10276
rect 41972 10220 41982 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 37436 10164 37492 10220
rect 2370 10108 2380 10164
rect 2436 10108 2446 10164
rect 5954 10108 5964 10164
rect 6020 10108 8540 10164
rect 8596 10108 8988 10164
rect 9044 10108 9054 10164
rect 10210 10108 10220 10164
rect 10276 10108 14252 10164
rect 14308 10108 14318 10164
rect 16818 10108 16828 10164
rect 16884 10108 17052 10164
rect 17108 10108 17118 10164
rect 17938 10108 17948 10164
rect 18004 10108 19292 10164
rect 19348 10108 19358 10164
rect 25666 10108 25676 10164
rect 25732 10108 26236 10164
rect 26292 10108 26302 10164
rect 29474 10108 29484 10164
rect 29540 10108 29708 10164
rect 29764 10108 29774 10164
rect 36082 10108 36092 10164
rect 36148 10108 36988 10164
rect 37044 10108 37436 10164
rect 37492 10108 37502 10164
rect 37650 10108 37660 10164
rect 37716 10108 41580 10164
rect 41636 10108 41646 10164
rect 2380 10052 2436 10108
rect 2380 9996 3276 10052
rect 3332 9996 3342 10052
rect 4946 9996 4956 10052
rect 5012 9996 7084 10052
rect 7140 9996 7150 10052
rect 7746 9996 7756 10052
rect 7812 9996 8988 10052
rect 9044 9996 9054 10052
rect 9762 9996 9772 10052
rect 9828 9996 13356 10052
rect 13412 9996 13422 10052
rect 14130 9996 14140 10052
rect 14196 9996 15596 10052
rect 15652 9996 15662 10052
rect 20850 9996 20860 10052
rect 20916 9996 21868 10052
rect 21924 9996 21934 10052
rect 22642 9996 22652 10052
rect 22708 9996 23772 10052
rect 23828 9996 24892 10052
rect 24948 9996 27580 10052
rect 27636 9996 27646 10052
rect 27794 9996 27804 10052
rect 27860 9996 30604 10052
rect 30660 9996 31724 10052
rect 31780 9996 31790 10052
rect 36204 9996 38780 10052
rect 38836 9996 40572 10052
rect 40628 9996 40638 10052
rect 2146 9884 2156 9940
rect 2212 9884 2716 9940
rect 2772 9884 2782 9940
rect 4162 9884 4172 9940
rect 4228 9884 4732 9940
rect 4788 9884 4798 9940
rect 6738 9884 6748 9940
rect 6804 9884 8092 9940
rect 8148 9884 8158 9940
rect 12786 9884 12796 9940
rect 12852 9884 12908 9940
rect 12964 9884 12974 9940
rect 14242 9884 14252 9940
rect 14308 9884 14924 9940
rect 14980 9884 16044 9940
rect 16100 9884 16110 9940
rect 17938 9884 17948 9940
rect 18004 9884 18620 9940
rect 18676 9884 18686 9940
rect 18946 9884 18956 9940
rect 19012 9884 19628 9940
rect 19684 9884 19694 9940
rect 21410 9884 21420 9940
rect 21476 9884 21980 9940
rect 22036 9884 22046 9940
rect 27458 9884 27468 9940
rect 27524 9884 28476 9940
rect 28532 9884 28542 9940
rect 33282 9884 33292 9940
rect 33348 9884 33740 9940
rect 33796 9884 33806 9940
rect 36204 9828 36260 9996
rect 37650 9884 37660 9940
rect 37716 9884 38668 9940
rect 38724 9884 38734 9940
rect 3042 9772 3052 9828
rect 3108 9772 3276 9828
rect 3332 9772 7644 9828
rect 7700 9772 7710 9828
rect 7970 9772 7980 9828
rect 8036 9772 9772 9828
rect 9828 9772 9838 9828
rect 12114 9772 12124 9828
rect 12180 9772 13692 9828
rect 13748 9772 13758 9828
rect 13906 9772 13916 9828
rect 13972 9772 15036 9828
rect 15092 9772 15102 9828
rect 15250 9772 15260 9828
rect 15316 9772 16492 9828
rect 16548 9772 16558 9828
rect 17714 9772 17724 9828
rect 17780 9772 19180 9828
rect 19236 9772 20860 9828
rect 20916 9772 21532 9828
rect 21588 9772 21598 9828
rect 22978 9772 22988 9828
rect 23044 9772 23548 9828
rect 23604 9772 26012 9828
rect 26068 9772 26460 9828
rect 26516 9772 26526 9828
rect 30034 9772 30044 9828
rect 30100 9772 31052 9828
rect 31108 9772 31388 9828
rect 31444 9772 31454 9828
rect 33842 9772 33852 9828
rect 33908 9772 34188 9828
rect 34244 9772 36204 9828
rect 36260 9772 36270 9828
rect 38098 9772 38108 9828
rect 38164 9772 38444 9828
rect 38500 9772 40124 9828
rect 40180 9772 41020 9828
rect 41076 9772 41086 9828
rect 1810 9660 1820 9716
rect 1876 9660 2156 9716
rect 2212 9660 2222 9716
rect 5394 9660 5404 9716
rect 5460 9660 9548 9716
rect 9604 9660 9614 9716
rect 10770 9660 10780 9716
rect 10836 9660 12684 9716
rect 12740 9660 12750 9716
rect 16790 9660 16828 9716
rect 16884 9660 16894 9716
rect 17826 9660 17836 9716
rect 17892 9660 19516 9716
rect 19572 9660 19582 9716
rect 19842 9660 19852 9716
rect 19908 9660 20412 9716
rect 20468 9660 20478 9716
rect 31154 9660 31164 9716
rect 31220 9660 35420 9716
rect 35476 9660 35644 9716
rect 35700 9660 36316 9716
rect 36372 9660 36382 9716
rect 38210 9660 38220 9716
rect 38276 9660 38780 9716
rect 38836 9660 38846 9716
rect 38994 9660 39004 9716
rect 39060 9660 39564 9716
rect 39620 9660 39630 9716
rect 5702 9548 5740 9604
rect 5796 9548 5806 9604
rect 6402 9548 6412 9604
rect 6468 9548 8204 9604
rect 8260 9548 8270 9604
rect 9958 9548 9996 9604
rect 10052 9548 10062 9604
rect 10854 9548 10892 9604
rect 10948 9548 10958 9604
rect 13010 9548 13020 9604
rect 13076 9548 18844 9604
rect 18900 9548 18910 9604
rect 19628 9548 19740 9604
rect 19796 9548 20300 9604
rect 20356 9548 20366 9604
rect 20514 9548 20524 9604
rect 20580 9548 21980 9604
rect 22036 9548 22046 9604
rect 33058 9548 33068 9604
rect 33124 9548 38556 9604
rect 38612 9548 41916 9604
rect 41972 9548 41982 9604
rect 19628 9492 19684 9548
rect 4162 9436 4172 9492
rect 4228 9436 6524 9492
rect 6580 9436 6590 9492
rect 7830 9436 7868 9492
rect 7924 9436 7934 9492
rect 8418 9436 8428 9492
rect 8484 9436 14588 9492
rect 14644 9436 14654 9492
rect 15138 9436 15148 9492
rect 15204 9436 19684 9492
rect 26338 9436 26348 9492
rect 26404 9436 27580 9492
rect 27636 9436 27646 9492
rect 30370 9436 30380 9492
rect 30436 9436 30940 9492
rect 30996 9436 31006 9492
rect 32022 9436 32060 9492
rect 32116 9436 32126 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4722 9324 4732 9380
rect 4788 9324 7196 9380
rect 7252 9324 7756 9380
rect 7812 9324 7822 9380
rect 12786 9324 12796 9380
rect 12852 9324 14700 9380
rect 14756 9324 19684 9380
rect 27682 9324 27692 9380
rect 27748 9324 32620 9380
rect 32676 9324 37436 9380
rect 37492 9324 38220 9380
rect 38276 9324 38286 9380
rect 19628 9268 19684 9324
rect 3266 9212 3276 9268
rect 3332 9212 6524 9268
rect 6580 9212 6590 9268
rect 7046 9212 7084 9268
rect 7140 9212 7150 9268
rect 13430 9212 13468 9268
rect 13524 9212 13534 9268
rect 16706 9212 16716 9268
rect 16772 9212 17836 9268
rect 17892 9212 17902 9268
rect 19628 9212 20636 9268
rect 20692 9212 21420 9268
rect 21476 9212 23436 9268
rect 23492 9212 23502 9268
rect 29810 9212 29820 9268
rect 29876 9212 33516 9268
rect 33572 9212 33582 9268
rect 34738 9212 34748 9268
rect 34804 9212 34814 9268
rect 6402 9100 6412 9156
rect 6468 9100 7532 9156
rect 7588 9100 7598 9156
rect 8978 9100 8988 9156
rect 9044 9100 12236 9156
rect 12292 9100 15316 9156
rect 4274 8988 4284 9044
rect 4340 8988 5852 9044
rect 5908 8988 5918 9044
rect 6262 8988 6300 9044
rect 6356 8988 6366 9044
rect 9874 8988 9884 9044
rect 9940 8988 10108 9044
rect 10164 8988 10174 9044
rect 15260 8932 15316 9100
rect 15484 9100 21084 9156
rect 21140 9100 21150 9156
rect 27682 9100 27692 9156
rect 27748 9100 30268 9156
rect 30324 9100 30334 9156
rect 15484 9044 15540 9100
rect 34748 9044 34804 9212
rect 35410 9100 35420 9156
rect 35476 9100 37548 9156
rect 37604 9100 37614 9156
rect 15474 8988 15484 9044
rect 15540 8988 15550 9044
rect 15810 8988 15820 9044
rect 15876 8988 16268 9044
rect 16324 8988 16334 9044
rect 16482 8988 16492 9044
rect 16548 8988 17612 9044
rect 17668 8988 17678 9044
rect 19842 8988 19852 9044
rect 19908 8988 21420 9044
rect 21476 8988 23660 9044
rect 23716 8988 23726 9044
rect 26002 8988 26012 9044
rect 26068 8988 28588 9044
rect 28644 8988 29596 9044
rect 29652 8988 31724 9044
rect 31780 8988 32508 9044
rect 32564 8988 32574 9044
rect 32946 8988 32956 9044
rect 33012 8988 33852 9044
rect 33908 8988 35644 9044
rect 35700 8988 36092 9044
rect 36148 8988 36158 9044
rect 38434 8988 38444 9044
rect 38500 8988 39676 9044
rect 39732 8988 40012 9044
rect 40068 8988 40078 9044
rect 5170 8876 5180 8932
rect 5236 8876 7084 8932
rect 7140 8876 8540 8932
rect 8596 8876 8606 8932
rect 10434 8876 10444 8932
rect 10500 8876 13580 8932
rect 13636 8876 13646 8932
rect 15260 8876 19180 8932
rect 19236 8876 19246 8932
rect 19404 8876 20860 8932
rect 20916 8876 25228 8932
rect 25284 8876 26236 8932
rect 26292 8876 26302 8932
rect 27794 8876 27804 8932
rect 27860 8876 30268 8932
rect 30324 8876 30334 8932
rect 31042 8876 31052 8932
rect 31108 8876 31836 8932
rect 31892 8876 31902 8932
rect 37538 8876 37548 8932
rect 37604 8876 39004 8932
rect 39060 8876 39070 8932
rect 19404 8820 19460 8876
rect 3938 8764 3948 8820
rect 4004 8764 8204 8820
rect 8260 8764 8270 8820
rect 8950 8764 8988 8820
rect 9044 8764 9054 8820
rect 9538 8764 9548 8820
rect 9604 8764 10780 8820
rect 10836 8764 10846 8820
rect 15110 8764 15148 8820
rect 15204 8764 18396 8820
rect 18452 8764 18462 8820
rect 19394 8764 19404 8820
rect 19460 8764 19470 8820
rect 24546 8764 24556 8820
rect 24612 8764 24892 8820
rect 24948 8764 24958 8820
rect 29138 8764 29148 8820
rect 29204 8764 30940 8820
rect 30996 8764 31006 8820
rect 36194 8764 36204 8820
rect 36260 8764 38668 8820
rect 38724 8764 38734 8820
rect 5282 8652 5292 8708
rect 5348 8652 10892 8708
rect 10948 8652 10958 8708
rect 11218 8652 11228 8708
rect 11284 8652 15876 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 15820 8596 15876 8652
rect 19404 8596 19460 8764
rect 30370 8652 30380 8708
rect 30436 8652 33628 8708
rect 33684 8652 33694 8708
rect 33954 8652 33964 8708
rect 34020 8652 34524 8708
rect 34580 8652 34590 8708
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 2146 8540 2156 8596
rect 2212 8540 3388 8596
rect 5926 8540 5964 8596
rect 6020 8540 6030 8596
rect 8204 8540 10444 8596
rect 10500 8540 10510 8596
rect 12898 8540 12908 8596
rect 12964 8540 13804 8596
rect 13860 8540 13870 8596
rect 15092 8540 15484 8596
rect 15540 8540 15550 8596
rect 15820 8540 19068 8596
rect 19124 8540 19460 8596
rect 21970 8540 21980 8596
rect 22036 8540 22764 8596
rect 22820 8540 22830 8596
rect 24210 8540 24220 8596
rect 24276 8540 32788 8596
rect 36082 8540 36092 8596
rect 36148 8540 37996 8596
rect 38052 8540 39340 8596
rect 39396 8540 39406 8596
rect 3332 8484 3388 8540
rect 8204 8484 8260 8540
rect 15092 8484 15148 8540
rect 32732 8484 32788 8540
rect 1922 8428 1932 8484
rect 1988 8428 2940 8484
rect 2996 8428 3006 8484
rect 3332 8428 6300 8484
rect 6356 8428 6366 8484
rect 6850 8428 6860 8484
rect 6916 8428 8204 8484
rect 8260 8428 8270 8484
rect 8530 8428 8540 8484
rect 8596 8428 8876 8484
rect 8932 8428 10332 8484
rect 10388 8428 15148 8484
rect 15810 8428 15820 8484
rect 15876 8428 16716 8484
rect 16772 8428 16782 8484
rect 20962 8428 20972 8484
rect 21028 8428 22204 8484
rect 22260 8428 22270 8484
rect 24882 8428 24892 8484
rect 24948 8428 27132 8484
rect 27188 8428 27198 8484
rect 32732 8428 40460 8484
rect 40516 8428 40526 8484
rect 40674 8428 40684 8484
rect 40740 8428 40750 8484
rect 40684 8372 40740 8428
rect 3042 8316 3052 8372
rect 3108 8316 8316 8372
rect 8372 8316 8382 8372
rect 13682 8316 13692 8372
rect 13748 8316 16996 8372
rect 19282 8316 19292 8372
rect 19348 8316 19852 8372
rect 19908 8316 19918 8372
rect 22418 8316 22428 8372
rect 22484 8316 26572 8372
rect 26628 8316 26638 8372
rect 28578 8316 28588 8372
rect 28644 8316 30044 8372
rect 30100 8316 30110 8372
rect 30716 8316 32060 8372
rect 32116 8316 32126 8372
rect 32498 8316 32508 8372
rect 32564 8316 34300 8372
rect 34356 8316 34366 8372
rect 39554 8316 39564 8372
rect 39620 8316 40124 8372
rect 40180 8316 40190 8372
rect 40684 8316 41244 8372
rect 41300 8316 41468 8372
rect 41524 8316 41534 8372
rect 2034 8204 2044 8260
rect 2100 8204 6300 8260
rect 6356 8204 6366 8260
rect 9986 8204 9996 8260
rect 10052 8204 11228 8260
rect 11284 8204 13132 8260
rect 13188 8204 13198 8260
rect 14130 8204 14140 8260
rect 14196 8204 15596 8260
rect 15652 8204 15662 8260
rect 16940 8148 16996 8316
rect 21410 8204 21420 8260
rect 21476 8204 26124 8260
rect 26180 8204 26190 8260
rect 26450 8204 26460 8260
rect 26516 8204 27804 8260
rect 27860 8204 28252 8260
rect 28308 8204 28318 8260
rect 29922 8204 29932 8260
rect 29988 8204 30492 8260
rect 30548 8204 30558 8260
rect 30716 8148 30772 8316
rect 40684 8260 40740 8316
rect 31378 8204 31388 8260
rect 31444 8204 32732 8260
rect 32788 8204 32798 8260
rect 33730 8204 33740 8260
rect 33796 8204 34748 8260
rect 34804 8204 35084 8260
rect 35140 8204 39228 8260
rect 39284 8204 40740 8260
rect 2258 8092 2268 8148
rect 2324 8092 3500 8148
rect 3556 8092 3566 8148
rect 5030 8092 5068 8148
rect 5124 8092 5134 8148
rect 13682 8092 13692 8148
rect 13748 8092 14812 8148
rect 14868 8092 14878 8148
rect 16930 8092 16940 8148
rect 16996 8092 18284 8148
rect 18340 8092 18350 8148
rect 19842 8092 19852 8148
rect 19908 8092 21868 8148
rect 21924 8092 21934 8148
rect 23874 8092 23884 8148
rect 23940 8092 30772 8148
rect 30930 8092 30940 8148
rect 30996 8092 33628 8148
rect 33684 8092 33964 8148
rect 34020 8092 41132 8148
rect 41188 8092 41198 8148
rect 1698 7980 1708 8036
rect 1764 7980 2380 8036
rect 2436 7980 3724 8036
rect 3780 7980 3790 8036
rect 4050 7980 4060 8036
rect 4116 7980 5628 8036
rect 5684 7980 5694 8036
rect 6626 7980 6636 8036
rect 6692 7980 7644 8036
rect 7700 7980 7710 8036
rect 8306 7980 8316 8036
rect 8372 7980 8764 8036
rect 8820 7980 8830 8036
rect 11554 7980 11564 8036
rect 11620 7980 14140 8036
rect 14196 7980 14206 8036
rect 19730 7980 19740 8036
rect 19796 7980 20300 8036
rect 20356 7980 21644 8036
rect 21700 7980 21710 8036
rect 30258 7980 30268 8036
rect 30324 7980 30604 8036
rect 30660 7980 30670 8036
rect 32050 7980 32060 8036
rect 32116 7980 32396 8036
rect 32452 7980 33740 8036
rect 33796 7980 33806 8036
rect 34066 7980 34076 8036
rect 34132 7980 36316 8036
rect 36372 7980 38220 8036
rect 38276 7980 38286 8036
rect 40674 7980 40684 8036
rect 40740 7980 41020 8036
rect 41076 7980 42028 8036
rect 42084 7980 42094 8036
rect 3378 7868 3388 7924
rect 3444 7868 3500 7924
rect 3556 7868 4844 7924
rect 4900 7868 10892 7924
rect 10948 7868 10958 7924
rect 13458 7868 13468 7924
rect 13524 7868 16044 7924
rect 16100 7868 16828 7924
rect 16884 7868 16894 7924
rect 25554 7868 25564 7924
rect 25620 7868 27020 7924
rect 27076 7868 27086 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 30604 7812 30660 7980
rect 31938 7868 31948 7924
rect 32004 7868 32732 7924
rect 32788 7868 35532 7924
rect 35588 7868 36204 7924
rect 36260 7868 36270 7924
rect 39778 7868 39788 7924
rect 39844 7868 40348 7924
rect 40404 7868 40414 7924
rect 2818 7756 2828 7812
rect 2884 7756 8428 7812
rect 8484 7756 8494 7812
rect 14466 7756 14476 7812
rect 14532 7756 15260 7812
rect 15316 7756 15326 7812
rect 17154 7756 17164 7812
rect 17220 7756 18620 7812
rect 18676 7756 18686 7812
rect 29810 7756 29820 7812
rect 29876 7756 30324 7812
rect 30604 7756 33964 7812
rect 34020 7756 34030 7812
rect 30268 7700 30324 7756
rect 6514 7644 6524 7700
rect 6580 7644 6860 7700
rect 6916 7644 6926 7700
rect 7298 7644 7308 7700
rect 7364 7644 8876 7700
rect 8932 7644 8942 7700
rect 9090 7644 9100 7700
rect 9156 7644 9884 7700
rect 9940 7644 9950 7700
rect 10742 7644 10780 7700
rect 10836 7644 10846 7700
rect 12674 7644 12684 7700
rect 12740 7644 15372 7700
rect 15428 7644 15438 7700
rect 16370 7644 16380 7700
rect 16436 7644 17724 7700
rect 17780 7644 17790 7700
rect 17910 7644 17948 7700
rect 18004 7644 18014 7700
rect 18274 7644 18284 7700
rect 18340 7644 20748 7700
rect 20804 7644 20814 7700
rect 22418 7644 22428 7700
rect 22484 7644 24444 7700
rect 24500 7644 24510 7700
rect 27570 7644 27580 7700
rect 27636 7644 29932 7700
rect 29988 7644 29998 7700
rect 30268 7644 33908 7700
rect 34290 7644 34300 7700
rect 34356 7644 36428 7700
rect 36484 7644 38332 7700
rect 38388 7644 38668 7700
rect 40226 7644 40236 7700
rect 40292 7644 40302 7700
rect 10780 7588 10836 7644
rect 33852 7588 33908 7644
rect 38612 7588 38668 7644
rect 2034 7532 2044 7588
rect 2100 7532 5740 7588
rect 5796 7532 6636 7588
rect 6692 7532 6702 7588
rect 7942 7532 7980 7588
rect 8036 7532 8046 7588
rect 8652 7532 12012 7588
rect 12068 7532 12078 7588
rect 25666 7532 25676 7588
rect 25732 7532 26460 7588
rect 26516 7532 26526 7588
rect 33842 7532 33852 7588
rect 33908 7532 33918 7588
rect 35522 7532 35532 7588
rect 35588 7532 37660 7588
rect 37716 7532 37726 7588
rect 38612 7532 39788 7588
rect 39844 7532 39854 7588
rect 8652 7476 8708 7532
rect 40236 7476 40292 7644
rect 1922 7420 1932 7476
rect 1988 7420 4732 7476
rect 4788 7420 4798 7476
rect 5506 7420 5516 7476
rect 5572 7420 5628 7476
rect 5684 7420 5694 7476
rect 6850 7420 6860 7476
rect 6916 7420 7308 7476
rect 7364 7420 8708 7476
rect 10518 7420 10556 7476
rect 10612 7420 10622 7476
rect 19618 7420 19628 7476
rect 19684 7420 19852 7476
rect 19908 7420 19918 7476
rect 20850 7420 20860 7476
rect 20916 7420 22092 7476
rect 22148 7420 22158 7476
rect 25778 7420 25788 7476
rect 25844 7420 26796 7476
rect 26852 7420 28476 7476
rect 28532 7420 28542 7476
rect 37660 7420 37884 7476
rect 37940 7420 38556 7476
rect 38612 7420 40292 7476
rect 5516 7364 5572 7420
rect 37660 7364 37716 7420
rect 4162 7308 4172 7364
rect 4228 7308 5572 7364
rect 5954 7308 5964 7364
rect 6020 7308 6748 7364
rect 6804 7308 6814 7364
rect 15586 7308 15596 7364
rect 15652 7308 19292 7364
rect 19348 7308 19358 7364
rect 19506 7308 19516 7364
rect 19572 7308 20188 7364
rect 20244 7308 20254 7364
rect 20514 7308 20524 7364
rect 20580 7308 21532 7364
rect 21588 7308 21598 7364
rect 23650 7308 23660 7364
rect 23716 7308 23884 7364
rect 23940 7308 23950 7364
rect 26226 7308 26236 7364
rect 26292 7308 26684 7364
rect 26740 7308 26750 7364
rect 30482 7308 30492 7364
rect 30548 7308 31276 7364
rect 31332 7308 31342 7364
rect 34860 7308 36876 7364
rect 36932 7308 36942 7364
rect 37650 7308 37660 7364
rect 37716 7308 37726 7364
rect 39666 7308 39676 7364
rect 39732 7308 41692 7364
rect 41748 7308 41758 7364
rect 34860 7252 34916 7308
rect 6626 7196 6636 7252
rect 6692 7196 7644 7252
rect 7700 7196 7710 7252
rect 8614 7196 8652 7252
rect 8708 7196 8718 7252
rect 9314 7196 9324 7252
rect 9380 7196 9996 7252
rect 10052 7196 10062 7252
rect 10994 7196 11004 7252
rect 11060 7196 27132 7252
rect 27188 7196 29820 7252
rect 29876 7196 32956 7252
rect 33012 7196 33022 7252
rect 34850 7196 34860 7252
rect 34916 7196 34926 7252
rect 35074 7196 35084 7252
rect 35140 7196 36316 7252
rect 36372 7196 40796 7252
rect 40852 7196 41580 7252
rect 41636 7196 41646 7252
rect 5926 7084 5964 7140
rect 6020 7084 6030 7140
rect 6290 7084 6300 7140
rect 6356 7084 6412 7140
rect 6468 7084 6478 7140
rect 7970 7084 7980 7140
rect 8036 7084 10556 7140
rect 10612 7084 10622 7140
rect 10882 7084 10892 7140
rect 10948 7084 17500 7140
rect 17556 7084 17566 7140
rect 26534 7084 26572 7140
rect 26628 7084 26638 7140
rect 28914 7084 28924 7140
rect 28980 7084 29652 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 29596 7028 29652 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 9314 6972 9324 7028
rect 9380 6972 19852 7028
rect 19908 6972 24556 7028
rect 24612 6972 24622 7028
rect 26786 6972 26796 7028
rect 26852 6972 29260 7028
rect 29316 6972 29326 7028
rect 29586 6972 29596 7028
rect 29652 6972 30828 7028
rect 30884 6972 32956 7028
rect 33012 6972 33022 7028
rect 33618 6972 33628 7028
rect 33684 6972 34188 7028
rect 34244 6972 34254 7028
rect 4610 6860 4620 6916
rect 4676 6860 8652 6916
rect 8708 6860 8718 6916
rect 9762 6860 9772 6916
rect 9828 6860 15148 6916
rect 15586 6860 15596 6916
rect 15652 6860 17052 6916
rect 17108 6860 19180 6916
rect 19236 6860 19246 6916
rect 23090 6860 23100 6916
rect 23156 6860 24332 6916
rect 24388 6860 26908 6916
rect 31154 6860 31164 6916
rect 31220 6860 34636 6916
rect 34692 6860 36652 6916
rect 36708 6860 38668 6916
rect 15092 6804 15148 6860
rect 3266 6748 3276 6804
rect 3332 6748 4284 6804
rect 4340 6748 4350 6804
rect 5058 6748 5068 6804
rect 5124 6748 6076 6804
rect 6132 6748 11228 6804
rect 11284 6748 11294 6804
rect 12338 6748 12348 6804
rect 12404 6748 13804 6804
rect 13860 6748 13870 6804
rect 15092 6748 16716 6804
rect 16772 6748 16782 6804
rect 18844 6692 18900 6860
rect 26852 6804 26908 6860
rect 38612 6804 38668 6860
rect 21746 6748 21756 6804
rect 21812 6748 25564 6804
rect 25620 6748 25630 6804
rect 26852 6748 28252 6804
rect 28308 6748 36764 6804
rect 36820 6748 36830 6804
rect 38612 6748 41020 6804
rect 41076 6748 41086 6804
rect 42354 6748 42364 6804
rect 42420 6748 42924 6804
rect 42980 6748 42990 6804
rect 4722 6636 4732 6692
rect 4788 6636 5068 6692
rect 5124 6636 5134 6692
rect 5618 6636 5628 6692
rect 5684 6636 5694 6692
rect 6850 6636 6860 6692
rect 6916 6636 13804 6692
rect 13860 6636 17388 6692
rect 17444 6636 17454 6692
rect 18834 6636 18844 6692
rect 18900 6636 18910 6692
rect 21746 6636 21756 6692
rect 21812 6636 21868 6692
rect 21924 6636 24220 6692
rect 24276 6636 24286 6692
rect 26198 6636 26236 6692
rect 26292 6636 26302 6692
rect 28690 6636 28700 6692
rect 28756 6636 30604 6692
rect 30660 6636 30670 6692
rect 34402 6636 34412 6692
rect 34468 6636 35980 6692
rect 36036 6636 36046 6692
rect 40114 6636 40124 6692
rect 40180 6636 41692 6692
rect 41748 6636 41758 6692
rect 5628 6580 5684 6636
rect 1474 6524 1484 6580
rect 1540 6524 2828 6580
rect 2884 6524 2894 6580
rect 5628 6524 7532 6580
rect 7588 6524 7598 6580
rect 10434 6524 10444 6580
rect 10500 6524 12460 6580
rect 12516 6524 12526 6580
rect 14130 6524 14140 6580
rect 14196 6524 14588 6580
rect 14644 6524 14654 6580
rect 15250 6524 15260 6580
rect 15316 6524 15354 6580
rect 18498 6524 18508 6580
rect 18564 6524 19292 6580
rect 19348 6524 19358 6580
rect 19516 6524 23884 6580
rect 23940 6524 23950 6580
rect 25666 6524 25676 6580
rect 25732 6524 30492 6580
rect 30548 6524 30558 6580
rect 19516 6468 19572 6524
rect 2706 6412 2716 6468
rect 2772 6412 5628 6468
rect 5684 6412 5694 6468
rect 9958 6412 9996 6468
rect 10052 6412 10062 6468
rect 12786 6412 12796 6468
rect 12852 6412 16940 6468
rect 16996 6412 17006 6468
rect 18386 6412 18396 6468
rect 18452 6412 19572 6468
rect 20626 6412 20636 6468
rect 20692 6412 24780 6468
rect 24836 6412 24846 6468
rect 27682 6412 27692 6468
rect 27748 6412 29820 6468
rect 29876 6412 29886 6468
rect 42018 6412 42028 6468
rect 42084 6412 42812 6468
rect 42868 6412 42878 6468
rect 13906 6300 13916 6356
rect 13972 6300 15372 6356
rect 15428 6300 17276 6356
rect 17332 6300 18620 6356
rect 18676 6300 19404 6356
rect 19460 6300 19470 6356
rect 21634 6300 21644 6356
rect 21700 6300 23996 6356
rect 24052 6300 24062 6356
rect 24210 6300 24220 6356
rect 24276 6300 25900 6356
rect 25956 6300 32732 6356
rect 32788 6300 33180 6356
rect 33236 6300 33246 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4162 6188 4172 6244
rect 4228 6188 7308 6244
rect 7364 6188 7374 6244
rect 8082 6188 8092 6244
rect 8148 6188 8876 6244
rect 8932 6188 11116 6244
rect 11172 6188 11182 6244
rect 14354 6188 14364 6244
rect 14420 6188 15708 6244
rect 15764 6188 16828 6244
rect 16884 6188 19068 6244
rect 19124 6188 19134 6244
rect 28914 6188 28924 6244
rect 28980 6188 29596 6244
rect 29652 6188 32844 6244
rect 32900 6188 32910 6244
rect 38612 6188 41916 6244
rect 41972 6188 41982 6244
rect 38612 6132 38668 6188
rect 9874 6076 9884 6132
rect 9940 6076 10108 6132
rect 10164 6076 10174 6132
rect 16930 6076 16940 6132
rect 16996 6076 20636 6132
rect 20692 6076 20702 6132
rect 24434 6076 24444 6132
rect 24500 6076 25676 6132
rect 25732 6076 25742 6132
rect 29362 6076 29372 6132
rect 29428 6076 31052 6132
rect 31108 6076 31118 6132
rect 31500 6076 32172 6132
rect 32228 6076 32238 6132
rect 33842 6076 33852 6132
rect 33908 6076 37660 6132
rect 37716 6076 38108 6132
rect 38164 6076 38668 6132
rect 40898 6076 40908 6132
rect 40964 6076 41804 6132
rect 41860 6076 41870 6132
rect 31500 6020 31556 6076
rect 1250 5964 1260 6020
rect 1316 5964 5068 6020
rect 5124 5964 5516 6020
rect 5572 5964 5582 6020
rect 6178 5964 6188 6020
rect 6244 5964 11564 6020
rect 11620 5964 15596 6020
rect 15652 5964 15662 6020
rect 15782 5964 15820 6020
rect 15876 5964 15886 6020
rect 16818 5964 16828 6020
rect 16884 5964 18396 6020
rect 18452 5964 18462 6020
rect 21746 5964 21756 6020
rect 21812 5964 22428 6020
rect 22484 5964 22494 6020
rect 28578 5964 28588 6020
rect 28644 5964 29036 6020
rect 29092 5964 29102 6020
rect 29922 5964 29932 6020
rect 29988 5964 31500 6020
rect 31556 5964 31566 6020
rect 31826 5964 31836 6020
rect 31892 5964 35868 6020
rect 35924 5964 35934 6020
rect 37538 5964 37548 6020
rect 37604 5964 39564 6020
rect 39620 5964 40348 6020
rect 40404 5964 40414 6020
rect 5170 5852 5180 5908
rect 5236 5852 13468 5908
rect 13524 5852 13534 5908
rect 17378 5852 17388 5908
rect 17444 5852 17724 5908
rect 17780 5852 21868 5908
rect 21924 5852 21934 5908
rect 22978 5852 22988 5908
rect 23044 5852 24220 5908
rect 24276 5852 24286 5908
rect 29810 5852 29820 5908
rect 29876 5852 30380 5908
rect 30436 5852 30446 5908
rect 32274 5852 32284 5908
rect 32340 5852 33740 5908
rect 33796 5852 33806 5908
rect 37426 5852 37436 5908
rect 37492 5852 38556 5908
rect 38612 5852 39340 5908
rect 39396 5852 39406 5908
rect 37436 5796 37492 5852
rect 6962 5740 6972 5796
rect 7028 5740 10220 5796
rect 10276 5740 10286 5796
rect 11442 5740 11452 5796
rect 11508 5740 13468 5796
rect 13524 5740 13534 5796
rect 32050 5740 32060 5796
rect 32116 5740 37492 5796
rect 9202 5628 9212 5684
rect 9268 5628 16828 5684
rect 16884 5628 16894 5684
rect 18508 5628 20300 5684
rect 20356 5628 24780 5684
rect 24836 5628 24846 5684
rect 32722 5628 32732 5684
rect 32788 5628 38332 5684
rect 38388 5628 38398 5684
rect 18508 5572 18564 5628
rect 18498 5516 18508 5572
rect 18564 5516 18574 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 5394 5404 5404 5460
rect 5460 5404 11900 5460
rect 11956 5404 11966 5460
rect 14214 5404 14252 5460
rect 14308 5404 14318 5460
rect 16706 5404 16716 5460
rect 16772 5404 21644 5460
rect 21700 5404 21710 5460
rect 5842 5292 5852 5348
rect 5908 5292 11004 5348
rect 11060 5292 11070 5348
rect 17042 5292 17052 5348
rect 17108 5292 20300 5348
rect 20356 5292 20366 5348
rect 24546 5292 24556 5348
rect 24612 5292 26460 5348
rect 26516 5292 26526 5348
rect 31378 5292 31388 5348
rect 31444 5292 33404 5348
rect 33460 5292 33470 5348
rect 34066 5292 34076 5348
rect 34132 5292 35980 5348
rect 36036 5292 36046 5348
rect 37874 5292 37884 5348
rect 37940 5292 38444 5348
rect 38500 5292 38510 5348
rect 38892 5292 41804 5348
rect 41860 5292 41870 5348
rect 38892 5236 38948 5292
rect 1810 5180 1820 5236
rect 1876 5180 3500 5236
rect 3556 5180 3566 5236
rect 4946 5180 4956 5236
rect 5012 5180 5628 5236
rect 5684 5180 5694 5236
rect 14802 5180 14812 5236
rect 14868 5180 16044 5236
rect 16100 5180 16110 5236
rect 24658 5180 24668 5236
rect 24724 5180 27804 5236
rect 27860 5180 27870 5236
rect 30706 5180 30716 5236
rect 30772 5180 31612 5236
rect 31668 5180 31678 5236
rect 32834 5180 32844 5236
rect 32900 5180 33628 5236
rect 33684 5180 33694 5236
rect 33954 5180 33964 5236
rect 34020 5180 38948 5236
rect 40114 5180 40124 5236
rect 40180 5180 41356 5236
rect 41412 5180 41422 5236
rect 1362 5068 1372 5124
rect 1428 5068 5852 5124
rect 5908 5068 6860 5124
rect 6916 5068 6926 5124
rect 7634 5068 7644 5124
rect 7700 5068 10108 5124
rect 10164 5068 10174 5124
rect 12562 5068 12572 5124
rect 12628 5068 18060 5124
rect 18116 5068 18126 5124
rect 19730 5068 19740 5124
rect 19796 5068 20524 5124
rect 20580 5068 20590 5124
rect 22194 5068 22204 5124
rect 22260 5068 22540 5124
rect 22596 5068 23212 5124
rect 23268 5068 23996 5124
rect 24052 5068 25788 5124
rect 25844 5068 25854 5124
rect 28690 5068 28700 5124
rect 28756 5068 29036 5124
rect 29092 5068 29932 5124
rect 29988 5068 31164 5124
rect 31220 5068 31230 5124
rect 31388 5068 32508 5124
rect 32564 5068 32574 5124
rect 35410 5068 35420 5124
rect 35476 5068 37884 5124
rect 37940 5068 37950 5124
rect 39442 5068 39452 5124
rect 39508 5068 40684 5124
rect 40740 5068 40750 5124
rect 19740 5012 19796 5068
rect 2482 4956 2492 5012
rect 2548 4956 3276 5012
rect 3332 4956 3342 5012
rect 4834 4956 4844 5012
rect 4900 4956 8428 5012
rect 8484 4956 8494 5012
rect 8978 4956 8988 5012
rect 9044 4956 12348 5012
rect 12404 4956 12414 5012
rect 17490 4956 17500 5012
rect 17556 4956 19796 5012
rect 20150 4956 20188 5012
rect 20244 4956 20254 5012
rect 22390 4956 22428 5012
rect 22484 4956 22494 5012
rect 26674 4956 26684 5012
rect 26740 4956 27468 5012
rect 27524 4956 27534 5012
rect 22428 4900 22484 4956
rect 31388 4900 31444 5068
rect 35074 4956 35084 5012
rect 35140 4956 41916 5012
rect 41972 4956 41982 5012
rect 1586 4844 1596 4900
rect 1652 4844 6636 4900
rect 6692 4844 7420 4900
rect 7476 4844 7486 4900
rect 14354 4844 14364 4900
rect 14420 4844 22092 4900
rect 22148 4844 22158 4900
rect 22428 4844 31444 4900
rect 4722 4732 4732 4788
rect 4788 4732 9884 4788
rect 9940 4732 15148 4788
rect 15204 4732 16716 4788
rect 16772 4732 16782 4788
rect 20514 4732 20524 4788
rect 20580 4732 23100 4788
rect 23156 4732 23166 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 6178 4620 6188 4676
rect 6244 4620 8988 4676
rect 9044 4620 9054 4676
rect 9762 4620 9772 4676
rect 9828 4620 10444 4676
rect 10500 4620 10510 4676
rect 14130 4620 14140 4676
rect 14196 4620 17612 4676
rect 17668 4620 17678 4676
rect 22306 4620 22316 4676
rect 22372 4620 42140 4676
rect 42196 4620 42206 4676
rect 2146 4508 2156 4564
rect 2212 4508 3388 4564
rect 6962 4508 6972 4564
rect 7028 4508 12012 4564
rect 12068 4508 12078 4564
rect 18274 4508 18284 4564
rect 18340 4508 22988 4564
rect 23044 4508 23054 4564
rect 23202 4508 23212 4564
rect 23268 4508 23884 4564
rect 23940 4508 23950 4564
rect 28466 4508 28476 4564
rect 28532 4508 32732 4564
rect 32788 4508 32798 4564
rect 40002 4508 40012 4564
rect 40068 4508 41244 4564
rect 41300 4508 41692 4564
rect 41748 4508 41758 4564
rect 3332 4452 3388 4508
rect 3332 4396 6524 4452
rect 6580 4396 6860 4452
rect 6916 4396 6926 4452
rect 7606 4396 7644 4452
rect 7700 4396 9212 4452
rect 9268 4396 9278 4452
rect 10546 4396 10556 4452
rect 10612 4396 11228 4452
rect 11284 4396 13916 4452
rect 13972 4396 16828 4452
rect 16884 4396 16894 4452
rect 21634 4396 21644 4452
rect 21700 4396 22204 4452
rect 22260 4396 22270 4452
rect 30818 4396 30828 4452
rect 30884 4396 33628 4452
rect 33684 4396 33694 4452
rect 39330 4396 39340 4452
rect 39396 4396 41580 4452
rect 41636 4396 41646 4452
rect 6860 4340 6916 4396
rect 6850 4284 6860 4340
rect 6916 4284 6926 4340
rect 12674 4284 12684 4340
rect 12740 4284 14700 4340
rect 14756 4284 14766 4340
rect 18134 4284 18172 4340
rect 18228 4284 18238 4340
rect 28802 4284 28812 4340
rect 28868 4284 31612 4340
rect 31668 4284 31678 4340
rect 31938 4284 31948 4340
rect 32004 4284 33852 4340
rect 33908 4284 33918 4340
rect 9090 4172 9100 4228
rect 9156 4172 10332 4228
rect 10388 4172 10398 4228
rect 28578 4172 28588 4228
rect 28644 4172 28700 4228
rect 28756 4172 28766 4228
rect 36082 4172 36092 4228
rect 36148 4172 38220 4228
rect 38276 4172 38286 4228
rect 4946 4060 4956 4116
rect 5012 4060 9996 4116
rect 10052 4060 10062 4116
rect 11218 4060 11228 4116
rect 11284 4060 21420 4116
rect 21476 4060 21486 4116
rect 38322 4060 38332 4116
rect 38388 4060 39900 4116
rect 39956 4060 39966 4116
rect 18722 3948 18732 4004
rect 18788 3948 19292 4004
rect 19348 3948 21532 4004
rect 21588 3948 21598 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 10658 3836 10668 3892
rect 10724 3836 11452 3892
rect 11508 3836 11518 3892
rect 21858 3836 21868 3892
rect 21924 3836 23548 3892
rect 23604 3836 24892 3892
rect 24948 3836 26908 3892
rect 39218 3836 39228 3892
rect 39284 3836 42812 3892
rect 42868 3836 42878 3892
rect 26852 3780 26908 3836
rect 3266 3724 3276 3780
rect 3332 3668 3388 3780
rect 6178 3724 6188 3780
rect 6244 3724 7868 3780
rect 7924 3724 7934 3780
rect 8866 3724 8876 3780
rect 8932 3724 10332 3780
rect 10388 3724 10556 3780
rect 10612 3724 10622 3780
rect 17714 3724 17724 3780
rect 17780 3724 22316 3780
rect 22372 3724 22382 3780
rect 26852 3724 40908 3780
rect 40964 3724 40974 3780
rect 3332 3612 6748 3668
rect 6804 3612 6814 3668
rect 12786 3612 12796 3668
rect 12852 3612 14028 3668
rect 14084 3612 14094 3668
rect 14578 3612 14588 3668
rect 14644 3612 15484 3668
rect 15540 3612 16492 3668
rect 16548 3612 16558 3668
rect 25330 3612 25340 3668
rect 25396 3612 27804 3668
rect 27860 3612 27870 3668
rect 28018 3612 28028 3668
rect 28084 3612 29932 3668
rect 29988 3612 29998 3668
rect 32162 3612 32172 3668
rect 32228 3612 33852 3668
rect 33908 3612 33918 3668
rect 39106 3612 39116 3668
rect 39172 3612 41468 3668
rect 41524 3612 41534 3668
rect 11666 3500 11676 3556
rect 11732 3500 13244 3556
rect 13300 3500 17164 3556
rect 17220 3500 17230 3556
rect 17602 3500 17612 3556
rect 17668 3500 18508 3556
rect 18564 3500 19516 3556
rect 19572 3500 19582 3556
rect 33394 3500 33404 3556
rect 33460 3500 35644 3556
rect 35700 3500 35710 3556
rect 40114 3500 40124 3556
rect 40180 3500 41580 3556
rect 41636 3500 41646 3556
rect 7858 3388 7868 3444
rect 7924 3388 11732 3444
rect 14690 3388 14700 3444
rect 14756 3388 15820 3444
rect 15876 3388 15886 3444
rect 21298 3388 21308 3444
rect 21364 3388 22540 3444
rect 22596 3388 23324 3444
rect 23380 3388 23390 3444
rect 23986 3388 23996 3444
rect 24052 3388 25452 3444
rect 25508 3388 25518 3444
rect 34738 3388 34748 3444
rect 34804 3388 37212 3444
rect 37268 3388 37278 3444
rect 37426 3388 37436 3444
rect 37492 3388 39004 3444
rect 39060 3388 39070 3444
rect 10556 3332 10612 3388
rect 11676 3332 11732 3388
rect 6374 3276 6412 3332
rect 6468 3276 6478 3332
rect 10546 3276 10556 3332
rect 10612 3276 10622 3332
rect 11676 3276 42588 3332
rect 42644 3276 42654 3332
rect 2818 3164 2828 3220
rect 2884 3164 7196 3220
rect 7252 3164 7262 3220
rect 15586 3164 15596 3220
rect 15652 3164 17724 3220
rect 17780 3164 17790 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 1026 3052 1036 3108
rect 1092 3052 10220 3108
rect 10276 3052 10286 3108
rect 4162 2940 4172 2996
rect 4228 2940 13916 2996
rect 13972 2940 13982 2996
rect 15922 2940 15932 2996
rect 15988 2940 42364 2996
rect 42420 2940 42430 2996
rect 16818 2828 16828 2884
rect 16884 2828 17276 2884
rect 17332 2828 42476 2884
rect 42532 2828 42542 2884
rect 7074 2716 7084 2772
rect 7140 2716 25788 2772
rect 25844 2716 25854 2772
rect 3826 2604 3836 2660
rect 3892 2604 42700 2660
rect 42756 2604 42766 2660
rect 1138 2492 1148 2548
rect 1204 2492 2268 2548
rect 2324 2492 42924 2548
rect 42980 2492 42990 2548
<< via3 >>
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 6860 25452 6916 25508
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 11116 24556 11172 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 23548 24108 23604 24164
rect 10780 23996 10836 24052
rect 4284 23660 4340 23716
rect 3836 23548 3892 23604
rect 7868 23548 7924 23604
rect 13804 23548 13860 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 9884 23212 9940 23268
rect 1820 22988 1876 23044
rect 2604 22988 2660 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 7420 22652 7476 22708
rect 10108 22540 10164 22596
rect 10892 22428 10948 22484
rect 10556 22316 10612 22372
rect 2156 22092 2212 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 6524 21868 6580 21924
rect 15820 21868 15876 21924
rect 1932 21756 1988 21812
rect 10108 21756 10164 21812
rect 11564 21756 11620 21812
rect 4844 21644 4900 21700
rect 3836 21532 3892 21588
rect 7420 21420 7476 21476
rect 18172 21420 18228 21476
rect 18620 21420 18676 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 6636 21084 6692 21140
rect 7532 20972 7588 21028
rect 14924 20972 14980 21028
rect 2604 20636 2660 20692
rect 8428 20636 8484 20692
rect 7980 20524 8036 20580
rect 12460 20524 12516 20580
rect 17948 20524 18004 20580
rect 3612 20412 3668 20468
rect 7196 20412 7252 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 7644 20300 7700 20356
rect 2268 20188 2324 20244
rect 16716 19852 16772 19908
rect 6748 19740 6804 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 6524 19516 6580 19572
rect 2156 19404 2212 19460
rect 5068 19404 5124 19460
rect 9212 19404 9268 19460
rect 13580 19404 13636 19460
rect 6524 19180 6580 19236
rect 16716 19180 16772 19236
rect 14924 19068 14980 19124
rect 8988 18956 9044 19012
rect 20188 18956 20244 19012
rect 5068 18844 5124 18900
rect 16828 18844 16884 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 7868 18620 7924 18676
rect 10444 18620 10500 18676
rect 4956 18508 5012 18564
rect 7532 18508 7588 18564
rect 12908 18508 12964 18564
rect 22876 18508 22932 18564
rect 1932 18396 1988 18452
rect 6524 18396 6580 18452
rect 8540 18396 8596 18452
rect 18508 18396 18564 18452
rect 2044 18284 2100 18340
rect 11564 18284 11620 18340
rect 12796 18284 12852 18340
rect 5404 18172 5460 18228
rect 7532 18172 7588 18228
rect 9884 18172 9940 18228
rect 20188 18172 20244 18228
rect 25228 18172 25284 18228
rect 3724 18060 3780 18116
rect 6412 18060 6468 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 8204 17836 8260 17892
rect 7420 17724 7476 17780
rect 23884 17724 23940 17780
rect 3276 17612 3332 17668
rect 6524 17612 6580 17668
rect 7196 17612 7252 17668
rect 7532 17612 7588 17668
rect 20188 17612 20244 17668
rect 2716 17500 2772 17556
rect 4172 17388 4228 17444
rect 5068 17388 5124 17444
rect 9212 17388 9268 17444
rect 13356 17388 13412 17444
rect 22092 17388 22148 17444
rect 22428 17388 22484 17444
rect 3164 17276 3220 17332
rect 4060 17276 4116 17332
rect 7980 17276 8036 17332
rect 15260 17276 15316 17332
rect 21756 17276 21812 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 6972 17164 7028 17220
rect 8428 17164 8484 17220
rect 8876 17164 8932 17220
rect 14028 17164 14084 17220
rect 18396 17164 18452 17220
rect 23660 17164 23716 17220
rect 2044 17052 2100 17108
rect 4956 17052 5012 17108
rect 22092 17052 22148 17108
rect 1932 16940 1988 16996
rect 2716 16940 2772 16996
rect 6300 16940 6356 16996
rect 13468 16940 13524 16996
rect 23996 16940 24052 16996
rect 7532 16828 7588 16884
rect 16268 16828 16324 16884
rect 16604 16828 16660 16884
rect 25228 16828 25284 16884
rect 3724 16716 3780 16772
rect 8652 16716 8708 16772
rect 15260 16716 15316 16772
rect 20524 16716 20580 16772
rect 7868 16604 7924 16660
rect 6860 16492 6916 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 5068 16380 5124 16436
rect 6972 16156 7028 16212
rect 8988 16156 9044 16212
rect 14028 15932 14084 15988
rect 2268 15820 2324 15876
rect 3164 15820 3220 15876
rect 4060 15820 4116 15876
rect 4956 15820 5012 15876
rect 18284 15820 18340 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 19180 15484 19236 15540
rect 19628 15484 19684 15540
rect 28700 15484 28756 15540
rect 3836 15372 3892 15428
rect 4060 15260 4116 15316
rect 22540 15260 22596 15316
rect 23324 15260 23380 15316
rect 27244 15148 27300 15204
rect 5068 14924 5124 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 3388 14812 3444 14868
rect 4284 14812 4340 14868
rect 7980 14700 8036 14756
rect 11676 14700 11732 14756
rect 15036 14700 15092 14756
rect 1932 14588 1988 14644
rect 5516 14588 5572 14644
rect 15932 14588 15988 14644
rect 7980 14476 8036 14532
rect 18396 14924 18452 14980
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 22876 14812 22932 14868
rect 21980 14588 22036 14644
rect 13356 14364 13412 14420
rect 3612 14252 3668 14308
rect 4060 14252 4116 14308
rect 4284 14252 4340 14308
rect 4956 14252 5012 14308
rect 6972 14252 7028 14308
rect 27580 14252 27636 14308
rect 3836 14140 3892 14196
rect 13580 14140 13636 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 16380 14028 16436 14084
rect 23100 14028 23156 14084
rect 8876 13916 8932 13972
rect 9996 13916 10052 13972
rect 5628 13692 5684 13748
rect 13580 13692 13636 13748
rect 3164 13580 3220 13636
rect 3724 13468 3780 13524
rect 10556 13468 10612 13524
rect 12796 13356 12852 13412
rect 15260 13356 15316 13412
rect 19628 13356 19684 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 14924 13244 14980 13300
rect 11676 13132 11732 13188
rect 6972 13020 7028 13076
rect 5068 12908 5124 12964
rect 5404 12908 5460 12964
rect 13356 12908 13412 12964
rect 8540 12796 8596 12852
rect 22540 12796 22596 12852
rect 10892 12684 10948 12740
rect 23100 12684 23156 12740
rect 26908 12572 26964 12628
rect 33628 12572 33684 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 18284 12460 18340 12516
rect 19180 12460 19236 12516
rect 22092 12460 22148 12516
rect 26796 12460 26852 12516
rect 4060 12348 4116 12404
rect 7084 12348 7140 12404
rect 7532 12348 7588 12404
rect 16380 12348 16436 12404
rect 4844 12236 4900 12292
rect 11564 12236 11620 12292
rect 15932 12236 15988 12292
rect 23660 12236 23716 12292
rect 24108 12124 24164 12180
rect 3836 12012 3892 12068
rect 21980 12012 22036 12068
rect 23324 12012 23380 12068
rect 26796 11900 26852 11956
rect 33628 11900 33684 11956
rect 27244 11788 27300 11844
rect 30380 11788 30436 11844
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 15036 11564 15092 11620
rect 23436 11564 23492 11620
rect 5068 11340 5124 11396
rect 5516 11340 5572 11396
rect 5740 11340 5796 11396
rect 6636 11340 6692 11396
rect 10108 11340 10164 11396
rect 12460 11340 12516 11396
rect 23436 11340 23492 11396
rect 29820 11340 29876 11396
rect 6524 11228 6580 11284
rect 9772 11116 9828 11172
rect 10108 11116 10164 11172
rect 25228 11116 25284 11172
rect 26796 11116 26852 11172
rect 1820 11004 1876 11060
rect 8204 11004 8260 11060
rect 13692 11004 13748 11060
rect 14252 11004 14308 11060
rect 15148 10892 15204 10948
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 24108 10780 24164 10836
rect 26908 10780 26964 10836
rect 11340 10668 11396 10724
rect 10332 10556 10388 10612
rect 18508 10556 18564 10612
rect 19180 10556 19236 10612
rect 37660 10892 37716 10948
rect 25228 10668 25284 10724
rect 26236 10668 26292 10724
rect 26796 10668 26852 10724
rect 38556 10332 38612 10388
rect 11340 10220 11396 10276
rect 23548 10220 23604 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 5964 10108 6020 10164
rect 37660 10108 37716 10164
rect 8988 9996 9044 10052
rect 9772 9996 9828 10052
rect 6748 9884 6804 9940
rect 12908 9884 12964 9940
rect 3276 9772 3332 9828
rect 16828 9660 16884 9716
rect 5740 9548 5796 9604
rect 9996 9548 10052 9604
rect 10892 9548 10948 9604
rect 7868 9436 7924 9492
rect 27580 9436 27636 9492
rect 32060 9436 32116 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 7084 9212 7140 9268
rect 13468 9212 13524 9268
rect 16716 9212 16772 9268
rect 8988 9100 9044 9156
rect 6300 8988 6356 9044
rect 9884 8988 9940 9044
rect 16268 8988 16324 9044
rect 19180 8876 19236 8932
rect 8988 8764 9044 8820
rect 15148 8764 15204 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 30380 8652 30436 8708
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 5964 8540 6020 8596
rect 6300 8428 6356 8484
rect 16716 8428 16772 8484
rect 26572 8316 26628 8372
rect 32060 8316 32116 8372
rect 5068 8092 5124 8148
rect 33628 8092 33684 8148
rect 32060 7980 32116 8036
rect 3388 7868 3444 7924
rect 10892 7868 10948 7924
rect 13468 7868 13524 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 18620 7756 18676 7812
rect 29820 7756 29876 7812
rect 10780 7644 10836 7700
rect 17948 7644 18004 7700
rect 5740 7532 5796 7588
rect 7980 7532 8036 7588
rect 5628 7420 5684 7476
rect 10556 7420 10612 7476
rect 15596 7308 15652 7364
rect 23884 7308 23940 7364
rect 6636 7196 6692 7252
rect 8652 7196 8708 7252
rect 5964 7084 6020 7140
rect 6300 7084 6356 7140
rect 10892 7084 10948 7140
rect 26572 7084 26628 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 8652 6860 8708 6916
rect 4284 6748 4340 6804
rect 13804 6748 13860 6804
rect 5068 6636 5124 6692
rect 21756 6636 21812 6692
rect 26236 6636 26292 6692
rect 28700 6636 28756 6692
rect 10444 6524 10500 6580
rect 15260 6524 15316 6580
rect 23884 6524 23940 6580
rect 9996 6412 10052 6468
rect 29820 6412 29876 6468
rect 23996 6300 24052 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 11116 6188 11172 6244
rect 10108 6076 10164 6132
rect 15596 5964 15652 6020
rect 15820 5964 15876 6020
rect 13468 5852 13524 5908
rect 38556 5852 38612 5908
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 14252 5404 14308 5460
rect 20524 5068 20580 5124
rect 20188 4956 20244 5012
rect 22428 4956 22484 5012
rect 20524 4732 20580 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 10444 4620 10500 4676
rect 23884 4508 23940 4564
rect 6860 4396 6916 4452
rect 7644 4396 7700 4452
rect 18172 4284 18228 4340
rect 28700 4172 28756 4228
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 10332 3724 10388 3780
rect 15820 3388 15876 3444
rect 6412 3276 6468 3332
rect 15596 3164 15652 3220
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 4172 2940 4228 2996
<< metal4 >>
rect 4448 40012 4768 40828
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 19808 40796 20128 40828
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4284 23716 4340 23726
rect 3836 23604 3892 23614
rect 1820 23044 1876 23054
rect 1820 11060 1876 22988
rect 2604 23044 2660 23054
rect 2156 22148 2212 22158
rect 1932 21812 1988 21822
rect 1932 18452 1988 21756
rect 2156 19460 2212 22092
rect 2604 20692 2660 22988
rect 2604 20626 2660 20636
rect 3836 21588 3892 23548
rect 3612 20468 3668 20478
rect 2156 19394 2212 19404
rect 2268 20244 2324 20254
rect 1932 18386 1988 18396
rect 2044 18340 2100 18350
rect 2044 17108 2100 18284
rect 2044 17042 2100 17052
rect 1932 16996 1988 17006
rect 1932 14644 1988 16940
rect 2268 15876 2324 20188
rect 3276 17668 3332 17678
rect 2716 17556 2772 17566
rect 2716 16996 2772 17500
rect 2716 16930 2772 16940
rect 3164 17332 3220 17342
rect 2268 15810 2324 15820
rect 3164 15876 3220 17276
rect 1932 14578 1988 14588
rect 3164 13636 3220 15820
rect 3164 13570 3220 13580
rect 1820 10994 1876 11004
rect 3276 9828 3332 17612
rect 3276 9762 3332 9772
rect 3388 14868 3444 14878
rect 3388 7924 3444 14812
rect 3612 14308 3668 20412
rect 3612 14242 3668 14252
rect 3724 18116 3780 18126
rect 3724 16772 3780 18060
rect 3724 13524 3780 16716
rect 3836 15428 3892 21532
rect 4172 17444 4228 17454
rect 4060 17332 4116 17342
rect 4060 15876 4116 17276
rect 4060 15810 4116 15820
rect 3836 15148 3892 15372
rect 4060 15316 4116 15326
rect 3836 15092 4004 15148
rect 3724 13458 3780 13468
rect 3836 14196 3892 14206
rect 3836 12068 3892 14140
rect 3948 12404 4004 15092
rect 4060 14308 4116 15260
rect 4060 14242 4116 14252
rect 4060 12404 4116 12414
rect 3948 12348 4060 12404
rect 4060 12338 4116 12348
rect 3836 12002 3892 12012
rect 3388 7858 3444 7868
rect 4172 2996 4228 17388
rect 4284 14868 4340 23660
rect 4284 14802 4340 14812
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 6860 25508 6916 25518
rect 6524 21924 6580 21934
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4284 14308 4340 14318
rect 4284 6804 4340 14252
rect 4284 6738 4340 6748
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4844 21700 4900 21710
rect 4844 12292 4900 21644
rect 6524 19572 6580 21868
rect 6524 19506 6580 19516
rect 6636 21140 6692 21150
rect 5068 19460 5124 19470
rect 5068 18900 5124 19404
rect 4956 18564 5012 18574
rect 4956 17108 5012 18508
rect 4956 17042 5012 17052
rect 5068 17444 5124 18844
rect 6524 19236 6580 19246
rect 6524 18452 6580 19180
rect 6524 18386 6580 18396
rect 5068 16436 5124 17388
rect 5068 16370 5124 16380
rect 5404 18228 5460 18238
rect 4956 15876 5012 15886
rect 4956 14308 5012 15820
rect 4956 14242 5012 14252
rect 5068 14980 5124 14990
rect 5068 12964 5124 14924
rect 5068 12898 5124 12908
rect 5404 12964 5460 18172
rect 6412 18116 6468 18126
rect 6300 16996 6356 17006
rect 5404 12898 5460 12908
rect 5516 14644 5572 14654
rect 4844 12226 4900 12236
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 5068 11396 5124 11406
rect 5068 8148 5124 11340
rect 5516 11396 5572 14588
rect 5516 11330 5572 11340
rect 5628 13748 5684 13758
rect 5068 6692 5124 8092
rect 5628 7476 5684 13692
rect 5740 11396 5796 11406
rect 5740 9604 5796 11340
rect 5740 7588 5796 9548
rect 5740 7522 5796 7532
rect 5964 10164 6020 10174
rect 5964 8596 6020 10108
rect 5628 7410 5684 7420
rect 5964 7140 6020 8540
rect 5964 7074 6020 7084
rect 6300 9044 6356 16940
rect 6300 8484 6356 8988
rect 6300 7140 6356 8428
rect 6300 7074 6356 7084
rect 5068 6626 5124 6636
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 6412 3332 6468 18060
rect 6524 17668 6580 17678
rect 6524 11284 6580 17612
rect 6524 11218 6580 11228
rect 6636 11396 6692 21084
rect 6636 7252 6692 11340
rect 6748 19796 6804 19806
rect 6748 9940 6804 19740
rect 6748 9874 6804 9884
rect 6860 16548 6916 25452
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 11116 24612 11172 24622
rect 10780 24052 10836 24062
rect 7868 23604 7924 23614
rect 7420 22708 7476 22718
rect 7420 21476 7476 22652
rect 7196 20468 7252 20478
rect 7196 17668 7252 20412
rect 7196 17602 7252 17612
rect 7420 17780 7476 21420
rect 7532 21028 7588 21038
rect 7532 18564 7588 20972
rect 7532 18498 7588 18508
rect 7644 20356 7700 20366
rect 6636 7186 6692 7196
rect 6860 4452 6916 16492
rect 6972 17220 7028 17230
rect 6972 16212 7028 17164
rect 7420 16884 7476 17724
rect 7532 18228 7588 18238
rect 7532 17668 7588 18172
rect 7532 17602 7588 17612
rect 7532 16884 7588 16894
rect 7420 16828 7532 16884
rect 6972 16146 7028 16156
rect 6972 14308 7028 14318
rect 6972 13076 7028 14252
rect 6972 13010 7028 13020
rect 7084 12404 7140 12414
rect 7084 9268 7140 12348
rect 7532 12404 7588 16828
rect 7532 12338 7588 12348
rect 7084 9202 7140 9212
rect 6860 4386 6916 4396
rect 7644 4452 7700 20300
rect 7868 18676 7924 23548
rect 9884 23268 9940 23278
rect 8428 20692 8484 20702
rect 7868 16660 7924 18620
rect 7868 9492 7924 16604
rect 7980 20580 8036 20590
rect 7980 17332 8036 20524
rect 7980 14756 8036 17276
rect 7980 14690 8036 14700
rect 8204 17892 8260 17902
rect 7868 9426 7924 9436
rect 7980 14532 8036 14542
rect 7980 7588 8036 14476
rect 8204 11060 8260 17836
rect 8428 17220 8484 20636
rect 9212 19460 9268 19470
rect 8988 19012 9044 19022
rect 8428 17154 8484 17164
rect 8540 18452 8596 18462
rect 8540 12852 8596 18396
rect 8876 17220 8932 17230
rect 8540 12786 8596 12796
rect 8652 16772 8708 16782
rect 8204 10994 8260 11004
rect 7980 7522 8036 7532
rect 8652 7252 8708 16716
rect 8876 13972 8932 17164
rect 8988 16212 9044 18956
rect 9212 17444 9268 19404
rect 9212 17378 9268 17388
rect 9884 18228 9940 23212
rect 8988 16146 9044 16156
rect 8876 13906 8932 13916
rect 9772 11172 9828 11182
rect 8988 10052 9044 10062
rect 8988 9156 9044 9996
rect 9772 10052 9828 11116
rect 9772 9986 9828 9996
rect 8988 8820 9044 9100
rect 9884 9044 9940 18172
rect 10108 22596 10164 22606
rect 10108 21812 10164 22540
rect 9884 8978 9940 8988
rect 9996 13972 10052 13982
rect 9996 9604 10052 13916
rect 10108 11396 10164 21756
rect 10556 22372 10612 22382
rect 10108 11330 10164 11340
rect 10444 18676 10500 18686
rect 8988 8754 9044 8764
rect 8652 6916 8708 7196
rect 8652 6850 8708 6860
rect 9996 6468 10052 9548
rect 9996 6402 10052 6412
rect 10108 11172 10164 11182
rect 10108 6132 10164 11116
rect 10108 6066 10164 6076
rect 10332 10612 10388 10622
rect 7644 4386 7700 4396
rect 10332 3780 10388 10556
rect 10444 6580 10500 18620
rect 10556 13524 10612 22316
rect 10556 7476 10612 13468
rect 10780 7700 10836 23996
rect 10892 22484 10948 22494
rect 10892 12740 10948 22428
rect 10892 9604 10948 12684
rect 10892 9538 10948 9548
rect 10780 7634 10836 7644
rect 10892 7924 10948 7934
rect 10556 7410 10612 7420
rect 10892 7140 10948 7868
rect 10892 7074 10948 7084
rect 10444 4676 10500 6524
rect 11116 6244 11172 24556
rect 13804 23604 13860 23614
rect 11564 21812 11620 21822
rect 11564 18340 11620 21756
rect 11564 12292 11620 18284
rect 12460 20580 12516 20590
rect 11676 14756 11732 14766
rect 11676 13188 11732 14700
rect 11676 13122 11732 13132
rect 11564 12226 11620 12236
rect 12460 11396 12516 20524
rect 13580 19460 13636 19470
rect 12908 18564 12964 18574
rect 12796 18340 12852 18350
rect 12796 13412 12852 18284
rect 12796 13346 12852 13356
rect 12460 11330 12516 11340
rect 11340 10724 11396 10734
rect 11340 10276 11396 10668
rect 11340 10210 11396 10220
rect 12908 9940 12964 18508
rect 13356 17444 13412 17454
rect 13356 14420 13412 17388
rect 13356 12964 13412 14364
rect 13356 12898 13412 12908
rect 13468 16996 13524 17006
rect 12908 9874 12964 9884
rect 13468 9268 13524 16940
rect 13580 15148 13636 19404
rect 13580 15092 13748 15148
rect 13580 14196 13636 14206
rect 13580 13748 13636 14140
rect 13580 13682 13636 13692
rect 13692 11060 13748 15092
rect 13692 10994 13748 11004
rect 13468 9202 13524 9212
rect 11116 6178 11172 6188
rect 13468 7924 13524 7934
rect 13468 5908 13524 7868
rect 13804 6804 13860 23548
rect 19808 23548 20128 25060
rect 35168 40012 35488 40828
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 15820 21924 15876 21934
rect 14924 21028 14980 21038
rect 14924 19124 14980 20972
rect 14028 17220 14084 17230
rect 14028 15988 14084 17164
rect 14028 15922 14084 15932
rect 14924 13300 14980 19068
rect 15260 17332 15316 17342
rect 15260 16772 15316 17276
rect 15260 16706 15316 16716
rect 14924 13234 14980 13244
rect 15036 14756 15092 14766
rect 15036 11620 15092 14700
rect 15036 11554 15092 11564
rect 15260 13412 15316 13422
rect 13804 6738 13860 6748
rect 14252 11060 14308 11070
rect 13468 5842 13524 5852
rect 14252 5460 14308 11004
rect 15148 10948 15204 10958
rect 15148 8820 15204 10892
rect 15148 8754 15204 8764
rect 15260 6580 15316 13356
rect 15260 6514 15316 6524
rect 15596 7364 15652 7374
rect 14252 5394 14308 5404
rect 15596 6020 15652 7308
rect 10444 4610 10500 4620
rect 10332 3714 10388 3724
rect 6412 3266 6468 3276
rect 15596 3220 15652 5964
rect 15820 6020 15876 21868
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 18172 21476 18228 21486
rect 17948 20580 18004 20590
rect 16716 19908 16772 19918
rect 16716 19236 16772 19852
rect 16268 16884 16324 16894
rect 15932 14644 15988 14654
rect 15932 12292 15988 14588
rect 15932 12226 15988 12236
rect 16268 9044 16324 16828
rect 16604 16884 16660 16894
rect 16604 15148 16660 16828
rect 16380 15092 16660 15148
rect 16380 14084 16436 15092
rect 16380 12404 16436 14028
rect 16380 12338 16436 12348
rect 16268 8978 16324 8988
rect 16716 9268 16772 19180
rect 16828 18900 16884 18910
rect 16828 9716 16884 18844
rect 16828 9650 16884 9660
rect 16716 8484 16772 9212
rect 16716 8418 16772 8428
rect 17948 7700 18004 20524
rect 17948 7634 18004 7644
rect 15820 3444 15876 5964
rect 18172 4340 18228 21420
rect 18620 21476 18676 21486
rect 18508 18452 18564 18462
rect 18396 17220 18452 17230
rect 18284 15876 18340 15886
rect 18284 12516 18340 15820
rect 18396 14980 18452 17164
rect 18396 14914 18452 14924
rect 18284 12450 18340 12460
rect 18508 10612 18564 18396
rect 18508 10546 18564 10556
rect 18620 7812 18676 21420
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 23548 24164 23604 24174
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 20188 19012 20244 19022
rect 20188 18228 20244 18956
rect 20188 18162 20244 18172
rect 22876 18564 22932 18574
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19180 15540 19236 15550
rect 19180 12516 19236 15484
rect 19628 15540 19684 15550
rect 19628 13412 19684 15484
rect 19628 13346 19684 13356
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19180 12450 19236 12460
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19180 10612 19236 10622
rect 19180 8932 19236 10556
rect 19180 8866 19236 8876
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 18620 7746 18676 7756
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 18172 4274 18228 4284
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 20188 17668 20244 17678
rect 20188 5012 20244 17612
rect 22092 17444 22148 17454
rect 21756 17332 21812 17342
rect 20188 4946 20244 4956
rect 20524 16772 20580 16782
rect 20524 5124 20580 16716
rect 21756 6692 21812 17276
rect 22092 17108 22148 17388
rect 21980 14644 22036 14654
rect 21980 12068 22036 14588
rect 22092 12516 22148 17052
rect 22092 12450 22148 12460
rect 22428 17444 22484 17454
rect 21980 12002 22036 12012
rect 21756 6626 21812 6636
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 20524 4788 20580 5068
rect 22428 5012 22484 17388
rect 22540 15316 22596 15326
rect 22540 12852 22596 15260
rect 22876 14868 22932 18508
rect 22876 14802 22932 14812
rect 23324 15316 23380 15326
rect 22540 12786 22596 12796
rect 23100 14084 23156 14094
rect 23100 12740 23156 14028
rect 23100 12674 23156 12684
rect 23324 12068 23380 15260
rect 23324 12002 23380 12012
rect 23436 11620 23492 11630
rect 23436 11396 23492 11564
rect 23436 11330 23492 11340
rect 23548 10276 23604 24108
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 25228 18228 25284 18238
rect 23884 17780 23940 17790
rect 23660 17220 23716 17230
rect 23660 12292 23716 17164
rect 23660 12226 23716 12236
rect 23548 10210 23604 10220
rect 22428 4946 22484 4956
rect 23884 7364 23940 17724
rect 23884 6580 23940 7308
rect 20524 4722 20580 4732
rect 15820 3378 15876 3388
rect 15596 3154 15652 3164
rect 19808 3164 20128 4676
rect 23884 4564 23940 6524
rect 23996 16996 24052 17006
rect 23996 6356 24052 16940
rect 25228 16884 25284 18172
rect 24108 12180 24164 12190
rect 24108 10836 24164 12124
rect 24108 10770 24164 10780
rect 25228 11172 25284 16828
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 28700 15540 28756 15550
rect 27244 15204 27300 15214
rect 26908 12628 26964 12638
rect 26796 12516 26852 12526
rect 26796 11956 26852 12460
rect 26796 11890 26852 11900
rect 25228 10724 25284 11116
rect 26796 11172 26852 11182
rect 25228 10658 25284 10668
rect 26236 10724 26292 10734
rect 26236 6692 26292 10668
rect 26796 10724 26852 11116
rect 26908 10836 26964 12572
rect 27244 11844 27300 15148
rect 27244 11778 27300 11788
rect 27580 14308 27636 14318
rect 26908 10770 26964 10780
rect 26796 10658 26852 10668
rect 27580 9492 27636 14252
rect 27580 9426 27636 9436
rect 26572 8372 26628 8382
rect 26572 7140 26628 8316
rect 26572 7074 26628 7084
rect 26236 6626 26292 6636
rect 28700 6692 28756 15484
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 33628 12628 33684 12638
rect 33628 11956 33684 12572
rect 30380 11844 30436 11854
rect 23996 6290 24052 6300
rect 23884 4498 23940 4508
rect 28700 4228 28756 6636
rect 29820 11396 29876 11406
rect 29820 7812 29876 11340
rect 30380 8708 30436 11788
rect 30380 8642 30436 8652
rect 32060 9492 32116 9502
rect 32060 8372 32116 9436
rect 32060 8036 32116 8316
rect 33628 8148 33684 11900
rect 33628 8082 33684 8092
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 37660 10948 37716 10958
rect 37660 10164 37716 10892
rect 37660 10098 37716 10108
rect 38556 10388 38612 10398
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 32060 7970 32116 7980
rect 29820 6468 29876 7756
rect 29820 6402 29876 6412
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 28700 4162 28756 4172
rect 35168 5516 35488 7028
rect 38556 5908 38612 10332
rect 38556 5842 38612 5852
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 4172 2930 4228 2940
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A1
timestamp 1669390400
transform -1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A2
timestamp 1669390400
transform -1 0 15008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1669390400
transform 1 0 40320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__A1
timestamp 1669390400
transform 1 0 24304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__A2
timestamp 1669390400
transform 1 0 40880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1669390400
transform -1 0 2016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A1
timestamp 1669390400
transform 1 0 19152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__I
timestamp 1669390400
transform 1 0 28000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A1
timestamp 1669390400
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A2
timestamp 1669390400
transform -1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__I
timestamp 1669390400
transform 1 0 26208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__I
timestamp 1669390400
transform 1 0 29792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A1
timestamp 1669390400
transform 1 0 41440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A2
timestamp 1669390400
transform -1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1669390400
transform 1 0 12320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1669390400
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A2
timestamp 1669390400
transform -1 0 27104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A1
timestamp 1669390400
transform 1 0 41552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A2
timestamp 1669390400
transform -1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1669390400
transform 1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A2
timestamp 1669390400
transform -1 0 34832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A1
timestamp 1669390400
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A2
timestamp 1669390400
transform -1 0 31696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A1
timestamp 1669390400
transform 1 0 35504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__A1
timestamp 1669390400
transform 1 0 40432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__A2
timestamp 1669390400
transform 1 0 39536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1669390400
transform 1 0 34832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A2
timestamp 1669390400
transform 1 0 40544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I
timestamp 1669390400
transform 1 0 41888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A1
timestamp 1669390400
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A2
timestamp 1669390400
transform 1 0 42000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A1
timestamp 1669390400
transform 1 0 41440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__A1
timestamp 1669390400
transform 1 0 41440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A1
timestamp 1669390400
transform 1 0 41664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A2
timestamp 1669390400
transform 1 0 41216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1669390400
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A1
timestamp 1669390400
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2
timestamp 1669390400
transform -1 0 5936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1669390400
transform 1 0 11760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1669390400
transform 1 0 6608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1669390400
transform 1 0 8064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1669390400
transform 1 0 2800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1669390400
transform -1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A2
timestamp 1669390400
transform -1 0 9632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__B
timestamp 1669390400
transform -1 0 10976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A1
timestamp 1669390400
transform 1 0 9072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1669390400
transform -1 0 11424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__B
timestamp 1669390400
transform -1 0 10192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A1
timestamp 1669390400
transform 1 0 20496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A2
timestamp 1669390400
transform -1 0 1904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__394__A4
timestamp 1669390400
transform 1 0 19600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A1
timestamp 1669390400
transform -1 0 3136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A2
timestamp 1669390400
transform -1 0 5152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1669390400
transform -1 0 18256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A1
timestamp 1669390400
transform -1 0 5152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1669390400
transform -1 0 13552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A3
timestamp 1669390400
transform 1 0 12208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A1
timestamp 1669390400
transform 1 0 9632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A2
timestamp 1669390400
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A2
timestamp 1669390400
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A3
timestamp 1669390400
transform 1 0 22848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__I
timestamp 1669390400
transform 1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__I
timestamp 1669390400
transform -1 0 7728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I
timestamp 1669390400
transform 1 0 14560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__I
timestamp 1669390400
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1669390400
transform 1 0 14672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1669390400
transform 1 0 15344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I
timestamp 1669390400
transform 1 0 23184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I
timestamp 1669390400
transform 1 0 20832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A2
timestamp 1669390400
transform -1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A1
timestamp 1669390400
transform 1 0 4704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A2
timestamp 1669390400
transform 1 0 3472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1669390400
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__415__I
timestamp 1669390400
transform 1 0 17584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A2
timestamp 1669390400
transform 1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1669390400
transform -1 0 5824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A2
timestamp 1669390400
transform 1 0 9632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__418__A3
timestamp 1669390400
transform -1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1669390400
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A2
timestamp 1669390400
transform 1 0 2016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__I
timestamp 1669390400
transform 1 0 22400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__I
timestamp 1669390400
transform 1 0 3584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1669390400
transform -1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1669390400
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__424__I
timestamp 1669390400
transform -1 0 1904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1669390400
transform -1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A1
timestamp 1669390400
transform -1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__426__A2
timestamp 1669390400
transform 1 0 9408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A1
timestamp 1669390400
transform 1 0 7616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A2
timestamp 1669390400
transform -1 0 7392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A3
timestamp 1669390400
transform -1 0 6944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A4
timestamp 1669390400
transform 1 0 8624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__428__I
timestamp 1669390400
transform -1 0 2576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__I
timestamp 1669390400
transform -1 0 7504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__B
timestamp 1669390400
transform -1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__A1
timestamp 1669390400
transform -1 0 26544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__431__A2
timestamp 1669390400
transform -1 0 26096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1669390400
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A2
timestamp 1669390400
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A1
timestamp 1669390400
transform 1 0 21504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A2
timestamp 1669390400
transform -1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__B
timestamp 1669390400
transform -1 0 22176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A1
timestamp 1669390400
transform 1 0 32816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A2
timestamp 1669390400
transform 1 0 33264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__A1
timestamp 1669390400
transform -1 0 21728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__A2
timestamp 1669390400
transform -1 0 23184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__B2
timestamp 1669390400
transform 1 0 24752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__438__I
timestamp 1669390400
transform 1 0 30688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A1
timestamp 1669390400
transform -1 0 25760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1669390400
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A1
timestamp 1669390400
transform 1 0 32032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A2
timestamp 1669390400
transform 1 0 28672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A2
timestamp 1669390400
transform -1 0 26208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__B2
timestamp 1669390400
transform 1 0 38304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A1
timestamp 1669390400
transform -1 0 29680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A2
timestamp 1669390400
transform 1 0 29904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A1
timestamp 1669390400
transform 1 0 28000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A2
timestamp 1669390400
transform -1 0 28672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A1
timestamp 1669390400
transform 1 0 31136 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__A2
timestamp 1669390400
transform -1 0 30464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__A1
timestamp 1669390400
transform -1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A2
timestamp 1669390400
transform 1 0 27664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__B
timestamp 1669390400
transform 1 0 27216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1669390400
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A2
timestamp 1669390400
transform 1 0 35392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1669390400
transform 1 0 10528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A1
timestamp 1669390400
transform 1 0 33936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A2
timestamp 1669390400
transform 1 0 33264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__A2
timestamp 1669390400
transform 1 0 33712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__A1
timestamp 1669390400
transform 1 0 36512 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A3
timestamp 1669390400
transform -1 0 29120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__A1
timestamp 1669390400
transform 1 0 34832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__B
timestamp 1669390400
transform 1 0 29792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__A1
timestamp 1669390400
transform 1 0 32144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A2
timestamp 1669390400
transform 1 0 33488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A1
timestamp 1669390400
transform -1 0 31024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__A2
timestamp 1669390400
transform 1 0 35952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A2
timestamp 1669390400
transform -1 0 34160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__B
timestamp 1669390400
transform 1 0 39760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1669390400
transform 1 0 40208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A1
timestamp 1669390400
transform 1 0 36064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A2
timestamp 1669390400
transform 1 0 38752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A1
timestamp 1669390400
transform -1 0 32144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A2
timestamp 1669390400
transform 1 0 32368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A3
timestamp 1669390400
transform 1 0 41104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__I
timestamp 1669390400
transform -1 0 31808 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A2
timestamp 1669390400
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__I
timestamp 1669390400
transform 1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A1
timestamp 1669390400
transform 1 0 41888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A2
timestamp 1669390400
transform 1 0 38864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__A2
timestamp 1669390400
transform -1 0 31808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__B
timestamp 1669390400
transform -1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A2
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1669390400
transform -1 0 35504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A3
timestamp 1669390400
transform -1 0 33936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__A2
timestamp 1669390400
transform 1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__A1
timestamp 1669390400
transform -1 0 35952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A1
timestamp 1669390400
transform 1 0 39648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A2
timestamp 1669390400
transform 1 0 36960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__A2
timestamp 1669390400
transform 1 0 39200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A1
timestamp 1669390400
transform 1 0 41888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A4
timestamp 1669390400
transform 1 0 37856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A2
timestamp 1669390400
transform 1 0 40992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__A2
timestamp 1669390400
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__A2
timestamp 1669390400
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A3
timestamp 1669390400
transform 1 0 37408 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A3
timestamp 1669390400
transform 1 0 39648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A3
timestamp 1669390400
transform 1 0 40096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A1
timestamp 1669390400
transform -1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__B
timestamp 1669390400
transform -1 0 9744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A1
timestamp 1669390400
transform -1 0 8288 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A2
timestamp 1669390400
transform -1 0 6496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1669390400
transform 1 0 7056 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A2
timestamp 1669390400
transform 1 0 8512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__I
timestamp 1669390400
transform 1 0 10976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A2
timestamp 1669390400
transform 1 0 10640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__B1
timestamp 1669390400
transform -1 0 8736 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__B2
timestamp 1669390400
transform 1 0 11200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A1
timestamp 1669390400
transform -1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A2
timestamp 1669390400
transform 1 0 5712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A1
timestamp 1669390400
transform 1 0 20048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A2
timestamp 1669390400
transform 1 0 20944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__B1
timestamp 1669390400
transform 1 0 19376 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__B2
timestamp 1669390400
transform 1 0 18928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__C
timestamp 1669390400
transform 1 0 21952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A2
timestamp 1669390400
transform -1 0 7504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__B1
timestamp 1669390400
transform -1 0 5824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__B2
timestamp 1669390400
transform -1 0 2800 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__C
timestamp 1669390400
transform -1 0 7056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1669390400
transform 1 0 2128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A2
timestamp 1669390400
transform -1 0 1904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A1
timestamp 1669390400
transform 1 0 2688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A2
timestamp 1669390400
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A1
timestamp 1669390400
transform 1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A2
timestamp 1669390400
transform 1 0 5264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__509__A2
timestamp 1669390400
transform 1 0 5600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A1
timestamp 1669390400
transform -1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A3
timestamp 1669390400
transform -1 0 6048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A2
timestamp 1669390400
transform -1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A3
timestamp 1669390400
transform 1 0 6384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__A2
timestamp 1669390400
transform 1 0 14000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__B1
timestamp 1669390400
transform -1 0 15120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__B2
timestamp 1669390400
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A1
timestamp 1669390400
transform 1 0 7168 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A2
timestamp 1669390400
transform 1 0 4816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1669390400
transform 1 0 3360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A2
timestamp 1669390400
transform 1 0 4368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A1
timestamp 1669390400
transform -1 0 3360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A2
timestamp 1669390400
transform -1 0 2352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A3
timestamp 1669390400
transform -1 0 2912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A1
timestamp 1669390400
transform 1 0 2352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A2
timestamp 1669390400
transform 1 0 3136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A1
timestamp 1669390400
transform -1 0 5152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A2
timestamp 1669390400
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A3
timestamp 1669390400
transform 1 0 3808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__A2
timestamp 1669390400
transform 1 0 8512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A2
timestamp 1669390400
transform 1 0 7728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__B1
timestamp 1669390400
transform -1 0 5600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__B2
timestamp 1669390400
transform -1 0 4256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__C
timestamp 1669390400
transform 1 0 6272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__B1
timestamp 1669390400
transform -1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__B2
timestamp 1669390400
transform -1 0 4592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A1
timestamp 1669390400
transform 1 0 3024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A2
timestamp 1669390400
transform -1 0 3696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__B
timestamp 1669390400
transform -1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A1
timestamp 1669390400
transform 1 0 7840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A2
timestamp 1669390400
transform -1 0 6944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A1
timestamp 1669390400
transform 1 0 3920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A2
timestamp 1669390400
transform 1 0 5936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1669390400
transform -1 0 1904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A1
timestamp 1669390400
transform 1 0 2576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A2
timestamp 1669390400
transform 1 0 2128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A1
timestamp 1669390400
transform -1 0 7840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A2
timestamp 1669390400
transform -1 0 7168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A1
timestamp 1669390400
transform 1 0 7952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A2
timestamp 1669390400
transform 1 0 6720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A2
timestamp 1669390400
transform 1 0 6496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A3
timestamp 1669390400
transform -1 0 6272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__B1
timestamp 1669390400
transform -1 0 4144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__B2
timestamp 1669390400
transform 1 0 4368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__C
timestamp 1669390400
transform 1 0 7392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__I
timestamp 1669390400
transform -1 0 2128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__B2
timestamp 1669390400
transform 1 0 3920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A1
timestamp 1669390400
transform -1 0 2800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A2
timestamp 1669390400
transform 1 0 3136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__I
timestamp 1669390400
transform -1 0 2688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__536__A2
timestamp 1669390400
transform 1 0 4256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1669390400
transform -1 0 4704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A2
timestamp 1669390400
transform -1 0 6160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__B
timestamp 1669390400
transform 1 0 7056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A1
timestamp 1669390400
transform -1 0 6384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A2
timestamp 1669390400
transform 1 0 6160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A1
timestamp 1669390400
transform -1 0 6832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B1
timestamp 1669390400
transform -1 0 5600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B2
timestamp 1669390400
transform 1 0 4368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__C
timestamp 1669390400
transform 1 0 6832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B2
timestamp 1669390400
transform 1 0 4816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A2
timestamp 1669390400
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__A1
timestamp 1669390400
transform 1 0 7504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__B
timestamp 1669390400
transform 1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A1
timestamp 1669390400
transform -1 0 2016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A2
timestamp 1669390400
transform 1 0 2688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1669390400
transform 1 0 4704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A2
timestamp 1669390400
transform 1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__A3
timestamp 1669390400
transform 1 0 7952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__A1
timestamp 1669390400
transform 1 0 10080 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__B1
timestamp 1669390400
transform -1 0 10192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__B2
timestamp 1669390400
transform 1 0 8512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__C
timestamp 1669390400
transform 1 0 9632 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__I
timestamp 1669390400
transform 1 0 2128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__B2
timestamp 1669390400
transform 1 0 7056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A1
timestamp 1669390400
transform -1 0 4704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A2
timestamp 1669390400
transform 1 0 3472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A1
timestamp 1669390400
transform -1 0 4144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A2
timestamp 1669390400
transform -1 0 1904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B1
timestamp 1669390400
transform -1 0 9632 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B2
timestamp 1669390400
transform 1 0 8960 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__C
timestamp 1669390400
transform -1 0 11088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__I
timestamp 1669390400
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B2
timestamp 1669390400
transform 1 0 8960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A1
timestamp 1669390400
transform -1 0 3248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A2
timestamp 1669390400
transform -1 0 2688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1669390400
transform 1 0 3920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__A1
timestamp 1669390400
transform -1 0 14784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__A2
timestamp 1669390400
transform -1 0 15232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A1
timestamp 1669390400
transform 1 0 10640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A2
timestamp 1669390400
transform 1 0 6944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A2
timestamp 1669390400
transform 1 0 11984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A1
timestamp 1669390400
transform -1 0 12544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__B1
timestamp 1669390400
transform -1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__B2
timestamp 1669390400
transform 1 0 10416 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__C
timestamp 1669390400
transform 1 0 11424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__B2
timestamp 1669390400
transform 1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A1
timestamp 1669390400
transform 1 0 10192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A2
timestamp 1669390400
transform 1 0 11312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__B
timestamp 1669390400
transform 1 0 14112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A1
timestamp 1669390400
transform -1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A2
timestamp 1669390400
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__B1
timestamp 1669390400
transform 1 0 14448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__C
timestamp 1669390400
transform -1 0 12992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A2
timestamp 1669390400
transform -1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__B2
timestamp 1669390400
transform 1 0 11648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A1
timestamp 1669390400
transform -1 0 7728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A1
timestamp 1669390400
transform -1 0 8624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A2
timestamp 1669390400
transform 1 0 8512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__596__A2
timestamp 1669390400
transform -1 0 6832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A2
timestamp 1669390400
transform 1 0 14000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A1
timestamp 1669390400
transform -1 0 13776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A2
timestamp 1669390400
transform -1 0 13104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__B1
timestamp 1669390400
transform 1 0 14896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__C
timestamp 1669390400
transform -1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__B1
timestamp 1669390400
transform 1 0 14448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__B2
timestamp 1669390400
transform 1 0 11872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1669390400
transform 1 0 14112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A2
timestamp 1669390400
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__A2
timestamp 1669390400
transform -1 0 13104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A2
timestamp 1669390400
transform -1 0 15680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A2
timestamp 1669390400
transform 1 0 15904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__A2
timestamp 1669390400
transform 1 0 16576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A1
timestamp 1669390400
transform 1 0 16912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A2
timestamp 1669390400
transform -1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__B1
timestamp 1669390400
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__C
timestamp 1669390400
transform -1 0 15456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__B1
timestamp 1669390400
transform 1 0 15008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__B2
timestamp 1669390400
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A1
timestamp 1669390400
transform 1 0 15568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A2
timestamp 1669390400
transform -1 0 12320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__A2
timestamp 1669390400
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__A3
timestamp 1669390400
transform 1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__616__I
timestamp 1669390400
transform -1 0 12096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__A1
timestamp 1669390400
transform 1 0 10416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__A2
timestamp 1669390400
transform 1 0 11200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A1
timestamp 1669390400
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A2
timestamp 1669390400
transform -1 0 11872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__A2
timestamp 1669390400
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__619__A3
timestamp 1669390400
transform -1 0 15904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__A1
timestamp 1669390400
transform -1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__620__A2
timestamp 1669390400
transform -1 0 6384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__A1
timestamp 1669390400
transform 1 0 16800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__621__A2
timestamp 1669390400
transform 1 0 16016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__A2
timestamp 1669390400
transform 1 0 14112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__A1
timestamp 1669390400
transform 1 0 18704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__A2
timestamp 1669390400
transform 1 0 16464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__B1
timestamp 1669390400
transform 1 0 16016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__C
timestamp 1669390400
transform -1 0 16240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__B1
timestamp 1669390400
transform -1 0 12544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__B2
timestamp 1669390400
transform -1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__625__I
timestamp 1669390400
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__626__A2
timestamp 1669390400
transform 1 0 17360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A1
timestamp 1669390400
transform -1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A2
timestamp 1669390400
transform -1 0 3248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A1
timestamp 1669390400
transform -1 0 6272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A2
timestamp 1669390400
transform -1 0 3360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__A1
timestamp 1669390400
transform -1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__629__A2
timestamp 1669390400
transform -1 0 16352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__630__A1
timestamp 1669390400
transform 1 0 10416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__630__A2
timestamp 1669390400
transform 1 0 9632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__A2
timestamp 1669390400
transform -1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__A3
timestamp 1669390400
transform 1 0 17360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__A1
timestamp 1669390400
transform 1 0 20272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__A2
timestamp 1669390400
transform 1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__B1
timestamp 1669390400
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__C
timestamp 1669390400
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__B1
timestamp 1669390400
transform -1 0 18032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__B2
timestamp 1669390400
transform 1 0 16576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A1
timestamp 1669390400
transform -1 0 16688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__A2
timestamp 1669390400
transform 1 0 16912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__A1
timestamp 1669390400
transform 1 0 16912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__636__A2
timestamp 1669390400
transform 1 0 15792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__637__I
timestamp 1669390400
transform -1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__A1
timestamp 1669390400
transform 1 0 24304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__639__A2
timestamp 1669390400
transform 1 0 31024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__A1
timestamp 1669390400
transform 1 0 23520 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__640__A2
timestamp 1669390400
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__641__A2
timestamp 1669390400
transform 1 0 23072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__A2
timestamp 1669390400
transform 1 0 7056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A1
timestamp 1669390400
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A2
timestamp 1669390400
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__B1
timestamp 1669390400
transform 1 0 18928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__C
timestamp 1669390400
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B1
timestamp 1669390400
transform -1 0 21168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B2
timestamp 1669390400
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__649__I
timestamp 1669390400
transform 1 0 30688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__A1
timestamp 1669390400
transform -1 0 10080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__A2
timestamp 1669390400
transform -1 0 8400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__A1
timestamp 1669390400
transform 1 0 11312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__652__I
timestamp 1669390400
transform 1 0 26768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__653__A2
timestamp 1669390400
transform -1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__A2
timestamp 1669390400
transform 1 0 14672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__654__A3
timestamp 1669390400
transform -1 0 20272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A3
timestamp 1669390400
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A1
timestamp 1669390400
transform -1 0 20720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A2
timestamp 1669390400
transform 1 0 18032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__B1
timestamp 1669390400
transform 1 0 18480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__C
timestamp 1669390400
transform 1 0 8288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A1
timestamp 1669390400
transform 1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A2
timestamp 1669390400
transform 1 0 32816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__659__A2
timestamp 1669390400
transform -1 0 19264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__A1
timestamp 1669390400
transform -1 0 13328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__A2
timestamp 1669390400
transform 1 0 18592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__A1
timestamp 1669390400
transform 1 0 19376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__A2
timestamp 1669390400
transform 1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A1
timestamp 1669390400
transform 1 0 18480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A2
timestamp 1669390400
transform 1 0 11648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__A3
timestamp 1669390400
transform 1 0 20944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A1
timestamp 1669390400
transform 1 0 18256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A2
timestamp 1669390400
transform -1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__B1
timestamp 1669390400
transform -1 0 17136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__B2
timestamp 1669390400
transform 1 0 20832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__B
timestamp 1669390400
transform 1 0 13664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__A1
timestamp 1669390400
transform -1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__A2
timestamp 1669390400
transform 1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__A2
timestamp 1669390400
transform -1 0 21504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A1
timestamp 1669390400
transform 1 0 21392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A2
timestamp 1669390400
transform 1 0 27888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__B2
timestamp 1669390400
transform 1 0 26656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__B
timestamp 1669390400
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A1
timestamp 1669390400
transform 1 0 25536 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A2
timestamp 1669390400
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__B
timestamp 1669390400
transform 1 0 21728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__A2
timestamp 1669390400
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__A2
timestamp 1669390400
transform 1 0 27104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__697__A2
timestamp 1669390400
transform -1 0 22960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__A1
timestamp 1669390400
transform 1 0 19824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__B2
timestamp 1669390400
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__B
timestamp 1669390400
transform -1 0 23856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A1
timestamp 1669390400
transform 1 0 27552 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__703__A2
timestamp 1669390400
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__A1
timestamp 1669390400
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1669390400
transform 1 0 36736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1669390400
transform 1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1669390400
transform 1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1669390400
transform -1 0 27552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1669390400
transform -1 0 29568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1669390400
transform 1 0 31136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1669390400
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1669390400
transform 1 0 33488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1669390400
transform 1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1669390400
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1669390400
transform 1 0 34272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1669390400
transform 1 0 36400 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1669390400
transform 1 0 42000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1669390400
transform 1 0 34384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1669390400
transform 1 0 35056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__CLK
timestamp 1669390400
transform 1 0 18256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__CLK
timestamp 1669390400
transform 1 0 2688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__CLK
timestamp 1669390400
transform -1 0 5152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__CLK
timestamp 1669390400
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1669390400
transform -1 0 3584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1669390400
transform 1 0 5600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1669390400
transform 1 0 10864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1669390400
transform 1 0 12432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1669390400
transform 1 0 13328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1669390400
transform 1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1669390400
transform 1 0 22400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__CLK
timestamp 1669390400
transform 1 0 16912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1669390400
transform 1 0 29008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__CLK
timestamp 1669390400
transform 1 0 28672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__CLK
timestamp 1669390400
transform -1 0 18256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__CLK
timestamp 1669390400
transform -1 0 26880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__741__CLK
timestamp 1669390400
transform 1 0 31808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__CLK
timestamp 1669390400
transform 1 0 29344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__CLK
timestamp 1669390400
transform 1 0 12320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__CLK
timestamp 1669390400
transform 1 0 13776 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__D
timestamp 1669390400
transform -1 0 16128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1669390400
transform -1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1669390400
transform 1 0 17584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1669390400
transform -1 0 24528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1669390400
transform 1 0 36736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform 1 0 21392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 15456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 17360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 20048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform 1 0 21504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform 1 0 21952 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 3024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 13552 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 4144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform -1 0 3808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform -1 0 3696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform 1 0 17808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 11984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform 1 0 18480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform -1 0 1904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 40544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1669390400
transform 1 0 27776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1669390400
transform -1 0 26992 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51
timestamp 1669390400
transform 1 0 7056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86
timestamp 1669390400
transform 1 0 10976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121
timestamp 1669390400
transform 1 0 14896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_149
timestamp 1669390400
transform 1 0 18032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_156
timestamp 1669390400
transform 1 0 18816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_195
timestamp 1669390400
transform 1 0 23184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_203
timestamp 1669390400
transform 1 0 24080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_207
timestamp 1669390400
transform 1 0 24528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_227
timestamp 1669390400
transform 1 0 26768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_243
timestamp 1669390400
transform 1 0 28560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_262
timestamp 1669390400
transform 1 0 30688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1669390400
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_297
timestamp 1669390400
transform 1 0 34608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1669390400
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_332
timestamp 1669390400
transform 1 0 38528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_348
timestamp 1669390400
transform 1 0 40320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_355
timestamp 1669390400
transform 1 0 41104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_357
timestamp 1669390400
transform 1 0 41328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_364
timestamp 1669390400
transform 1 0 42112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_9
timestamp 1669390400
transform 1 0 2352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_13
timestamp 1669390400
transform 1 0 2800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_43
timestamp 1669390400
transform 1 0 6160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_52
timestamp 1669390400
transform 1 0 7168 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1669390400
transform 1 0 10080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_109
timestamp 1669390400
transform 1 0 13552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_140
timestamp 1669390400
transform 1 0 17024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_158
timestamp 1669390400
transform 1 0 19040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_160
timestamp 1669390400
transform 1 0 19264 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_190
timestamp 1669390400
transform 1 0 22624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_206
timestamp 1669390400
transform 1 0 24416 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_245
timestamp 1669390400
transform 1 0 28784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_249
timestamp 1669390400
transform 1 0 29232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_265
timestamp 1669390400
transform 1 0 31024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_275
timestamp 1669390400
transform 1 0 32144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_293
timestamp 1669390400
transform 1 0 34160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_295
timestamp 1669390400
transform 1 0 34384 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_325
timestamp 1669390400
transform 1 0 37744 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_341
timestamp 1669390400
transform 1 0 39536 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_349
timestamp 1669390400
transform 1 0 40432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_353
timestamp 1669390400
transform 1 0 40880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_364
timestamp 1669390400
transform 1 0 42112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_5
timestamp 1669390400
transform 1 0 1904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_16
timestamp 1669390400
transform 1 0 3136 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_42
timestamp 1669390400
transform 1 0 6048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_60
timestamp 1669390400
transform 1 0 8064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_91
timestamp 1669390400
transform 1 0 11536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_102
timestamp 1669390400
transform 1 0 12768 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_117
timestamp 1669390400
transform 1 0 14448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_135
timestamp 1669390400
transform 1 0 16464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_166
timestamp 1669390400
transform 1 0 19936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_181
timestamp 1669390400
transform 1 0 21616 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_191
timestamp 1669390400
transform 1 0 22736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_198
timestamp 1669390400
transform 1 0 23520 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_229
timestamp 1669390400
transform 1 0 26992 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_245
timestamp 1669390400
transform 1 0 28784 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_283
timestamp 1669390400
transform 1 0 33040 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_293
timestamp 1669390400
transform 1 0 34160 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_297
timestamp 1669390400
transform 1 0 34608 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_306
timestamp 1669390400
transform 1 0 35616 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_328
timestamp 1669390400
transform 1 0 38080 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_332
timestamp 1669390400
transform 1 0 38528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_348
timestamp 1669390400
transform 1 0 40320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_32
timestamp 1669390400
transform 1 0 4928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_34
timestamp 1669390400
transform 1 0 5152 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_51
timestamp 1669390400
transform 1 0 7056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_53
timestamp 1669390400
transform 1 0 7280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_83
timestamp 1669390400
transform 1 0 10640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_93
timestamp 1669390400
transform 1 0 11760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_111
timestamp 1669390400
transform 1 0 13776 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_117
timestamp 1669390400
transform 1 0 14448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_135
timestamp 1669390400
transform 1 0 16464 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_148
timestamp 1669390400
transform 1 0 17920 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_166
timestamp 1669390400
transform 1 0 19936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_197
timestamp 1669390400
transform 1 0 23408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_201
timestamp 1669390400
transform 1 0 23856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_218
timestamp 1669390400
transform 1 0 25760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_220
timestamp 1669390400
transform 1 0 25984 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_229
timestamp 1669390400
transform 1 0 26992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_239
timestamp 1669390400
transform 1 0 28112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_245
timestamp 1669390400
transform 1 0 28784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_256
timestamp 1669390400
transform 1 0 30016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_266
timestamp 1669390400
transform 1 0 31136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_276
timestamp 1669390400
transform 1 0 32256 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_294
timestamp 1669390400
transform 1 0 34272 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_325
timestamp 1669390400
transform 1 0 37744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_343
timestamp 1669390400
transform 1 0 39760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_351
timestamp 1669390400
transform 1 0 40656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_364
timestamp 1669390400
transform 1 0 42112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_9
timestamp 1669390400
transform 1 0 2352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_27
timestamp 1669390400
transform 1 0 4368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_49
timestamp 1669390400
transform 1 0 6832 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_53
timestamp 1669390400
transform 1 0 7280 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_67
timestamp 1669390400
transform 1 0 8848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_74
timestamp 1669390400
transform 1 0 9632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_84
timestamp 1669390400
transform 1 0 10752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_94
timestamp 1669390400
transform 1 0 11872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_118
timestamp 1669390400
transform 1 0 14560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_133
timestamp 1669390400
transform 1 0 16240 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_146
timestamp 1669390400
transform 1 0 17696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_150
timestamp 1669390400
transform 1 0 18144 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_162
timestamp 1669390400
transform 1 0 19488 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_166
timestamp 1669390400
transform 1 0 19936 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_188
timestamp 1669390400
transform 1 0 22400 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_242
timestamp 1669390400
transform 1 0 28448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1669390400
transform 1 0 28896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_257
timestamp 1669390400
transform 1 0 30128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_263
timestamp 1669390400
transform 1 0 30800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_294
timestamp 1669390400
transform 1 0 34272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_306
timestamp 1669390400
transform 1 0 35616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_331
timestamp 1669390400
transform 1 0 38416 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_333
timestamp 1669390400
transform 1 0 38640 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_348
timestamp 1669390400
transform 1 0 40320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_358
timestamp 1669390400
transform 1 0 41440 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_360
timestamp 1669390400
transform 1 0 41664 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_365
timestamp 1669390400
transform 1 0 42224 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_32
timestamp 1669390400
transform 1 0 4928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_34
timestamp 1669390400
transform 1 0 5152 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_45
timestamp 1669390400
transform 1 0 6384 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_47
timestamp 1669390400
transform 1 0 6608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_56
timestamp 1669390400
transform 1 0 7616 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_76
timestamp 1669390400
transform 1 0 9856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_88
timestamp 1669390400
transform 1 0 11200 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_140
timestamp 1669390400
transform 1 0 17024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_152
timestamp 1669390400
transform 1 0 18368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_165
timestamp 1669390400
transform 1 0 19824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_167
timestamp 1669390400
transform 1 0 20048 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_170
timestamp 1669390400
transform 1 0 20384 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_201
timestamp 1669390400
transform 1 0 23856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_209
timestamp 1669390400
transform 1 0 24752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_222
timestamp 1669390400
transform 1 0 26208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_228
timestamp 1669390400
transform 1 0 26880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_238
timestamp 1669390400
transform 1 0 28000 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_269
timestamp 1669390400
transform 1 0 31472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_271
timestamp 1669390400
transform 1 0 31696 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_280
timestamp 1669390400
transform 1 0 32704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_293
timestamp 1669390400
transform 1 0 34160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_326
timestamp 1669390400
transform 1 0 37856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_332
timestamp 1669390400
transform 1 0 38528 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_348
timestamp 1669390400
transform 1 0 40320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_364
timestamp 1669390400
transform 1 0 42112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_7
timestamp 1669390400
transform 1 0 2128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_16
timestamp 1669390400
transform 1 0 3136 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_27
timestamp 1669390400
transform 1 0 4368 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_49
timestamp 1669390400
transform 1 0 6832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_53
timestamp 1669390400
transform 1 0 7280 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_63
timestamp 1669390400
transform 1 0 8400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_73
timestamp 1669390400
transform 1 0 9520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_104
timestamp 1669390400
transform 1 0 12992 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_120
timestamp 1669390400
transform 1 0 14784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_126
timestamp 1669390400
transform 1 0 15456 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_136
timestamp 1669390400
transform 1 0 16576 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_147
timestamp 1669390400
transform 1 0 17808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_153
timestamp 1669390400
transform 1 0 18480 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_166
timestamp 1669390400
transform 1 0 19936 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_168
timestamp 1669390400
transform 1 0 20160 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_181
timestamp 1669390400
transform 1 0 21616 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_190
timestamp 1669390400
transform 1 0 22624 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1669390400
transform 1 0 28448 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_246
timestamp 1669390400
transform 1 0 28896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_262
timestamp 1669390400
transform 1 0 30688 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_270
timestamp 1669390400
transform 1 0 31584 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_274
timestamp 1669390400
transform 1 0 32032 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_276
timestamp 1669390400
transform 1 0 32256 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_285
timestamp 1669390400
transform 1 0 33264 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_293
timestamp 1669390400
transform 1 0 34160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_301
timestamp 1669390400
transform 1 0 35056 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_308
timestamp 1669390400
transform 1 0 35840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_315
timestamp 1669390400
transform 1 0 36624 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_328
timestamp 1669390400
transform 1 0 38080 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_335
timestamp 1669390400
transform 1 0 38864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_343
timestamp 1669390400
transform 1 0 39760 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_349
timestamp 1669390400
transform 1 0 40432 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_353
timestamp 1669390400
transform 1 0 40880 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_357
timestamp 1669390400
transform 1 0 41328 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_361
timestamp 1669390400
transform 1 0 41776 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_365
timestamp 1669390400
transform 1 0 42224 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_32
timestamp 1669390400
transform 1 0 4928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1669390400
transform 1 0 5600 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_48
timestamp 1669390400
transform 1 0 6720 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_58
timestamp 1669390400
transform 1 0 7840 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_60
timestamp 1669390400
transform 1 0 8064 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1669390400
transform 1 0 8960 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_83
timestamp 1669390400
transform 1 0 10640 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_85
timestamp 1669390400
transform 1 0 10864 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_94
timestamp 1669390400
transform 1 0 11872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_104
timestamp 1669390400
transform 1 0 12992 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_117
timestamp 1669390400
transform 1 0 14448 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_121
timestamp 1669390400
transform 1 0 14896 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_130
timestamp 1669390400
transform 1 0 15904 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_139
timestamp 1669390400
transform 1 0 16912 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_153
timestamp 1669390400
transform 1 0 18480 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_163
timestamp 1669390400
transform 1 0 19600 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_167
timestamp 1669390400
transform 1 0 20048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_176
timestamp 1669390400
transform 1 0 21056 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_178
timestamp 1669390400
transform 1 0 21280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_181
timestamp 1669390400
transform 1 0 21616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_245
timestamp 1669390400
transform 1 0 28784 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_253
timestamp 1669390400
transform 1 0 29680 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_261
timestamp 1669390400
transform 1 0 30576 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_269
timestamp 1669390400
transform 1 0 31472 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_277
timestamp 1669390400
transform 1 0 32368 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_281
timestamp 1669390400
transform 1 0 32816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_292
timestamp 1669390400
transform 1 0 34048 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_325
timestamp 1669390400
transform 1 0 37744 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_335
timestamp 1669390400
transform 1 0 38864 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_341
timestamp 1669390400
transform 1 0 39536 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_345
timestamp 1669390400
transform 1 0 39984 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_349
timestamp 1669390400
transform 1 0 40432 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_353
timestamp 1669390400
transform 1 0 40880 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_360
timestamp 1669390400
transform 1 0 41664 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_364
timestamp 1669390400
transform 1 0 42112 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_9
timestamp 1669390400
transform 1 0 2352 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_17
timestamp 1669390400
transform 1 0 3248 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_28
timestamp 1669390400
transform 1 0 4480 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_49
timestamp 1669390400
transform 1 0 6832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_51
timestamp 1669390400
transform 1 0 7056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_60
timestamp 1669390400
transform 1 0 8064 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_70
timestamp 1669390400
transform 1 0 9184 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1669390400
transform 1 0 10416 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_88
timestamp 1669390400
transform 1 0 11200 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_98
timestamp 1669390400
transform 1 0 12320 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_118
timestamp 1669390400
transform 1 0 14560 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_126
timestamp 1669390400
transform 1 0 15456 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_128
timestamp 1669390400
transform 1 0 15680 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_135
timestamp 1669390400
transform 1 0 16464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_143
timestamp 1669390400
transform 1 0 17360 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_149
timestamp 1669390400
transform 1 0 18032 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_159
timestamp 1669390400
transform 1 0 19152 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_166
timestamp 1669390400
transform 1 0 19936 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_189
timestamp 1669390400
transform 1 0 22512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_193
timestamp 1669390400
transform 1 0 22960 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_224
timestamp 1669390400
transform 1 0 26432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_228
timestamp 1669390400
transform 1 0 26880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_230
timestamp 1669390400
transform 1 0 27104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_239
timestamp 1669390400
transform 1 0 28112 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_260
timestamp 1669390400
transform 1 0 30464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_275
timestamp 1669390400
transform 1 0 32144 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_306
timestamp 1669390400
transform 1 0 35616 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_313
timestamp 1669390400
transform 1 0 36400 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1669390400
transform 1 0 36848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_330
timestamp 1669390400
transform 1 0 38304 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_338
timestamp 1669390400
transform 1 0 39200 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_344
timestamp 1669390400
transform 1 0 39872 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_348
timestamp 1669390400
transform 1 0 40320 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_352
timestamp 1669390400
transform 1 0 40768 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_356
timestamp 1669390400
transform 1 0 41216 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_360
timestamp 1669390400
transform 1 0 41664 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_364
timestamp 1669390400
transform 1 0 42112 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_19
timestamp 1669390400
transform 1 0 3472 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_21
timestamp 1669390400
transform 1 0 3696 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_31
timestamp 1669390400
transform 1 0 4816 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_40
timestamp 1669390400
transform 1 0 5824 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_49
timestamp 1669390400
transform 1 0 6832 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_59
timestamp 1669390400
transform 1 0 7952 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_61
timestamp 1669390400
transform 1 0 8176 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_85
timestamp 1669390400
transform 1 0 10864 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_91
timestamp 1669390400
transform 1 0 11536 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_122
timestamp 1669390400
transform 1 0 15008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_129
timestamp 1669390400
transform 1 0 15792 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_150
timestamp 1669390400
transform 1 0 18144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_202
timestamp 1669390400
transform 1 0 23968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_248
timestamp 1669390400
transform 1 0 29120 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_295
timestamp 1669390400
transform 1 0 34384 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_302
timestamp 1669390400
transform 1 0 35168 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_306
timestamp 1669390400
transform 1 0 35616 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_313
timestamp 1669390400
transform 1 0 36400 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_320
timestamp 1669390400
transform 1 0 37184 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_324
timestamp 1669390400
transform 1 0 37632 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_332
timestamp 1669390400
transform 1 0 38528 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_336
timestamp 1669390400
transform 1 0 38976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_340
timestamp 1669390400
transform 1 0 39424 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_344
timestamp 1669390400
transform 1 0 39872 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_348
timestamp 1669390400
transform 1 0 40320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_352
timestamp 1669390400
transform 1 0 40768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_360
timestamp 1669390400
transform 1 0 41664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_364
timestamp 1669390400
transform 1 0 42112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_32
timestamp 1669390400
transform 1 0 4928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_49
timestamp 1669390400
transform 1 0 6832 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_59
timestamp 1669390400
transform 1 0 7952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_61
timestamp 1669390400
transform 1 0 8176 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_64
timestamp 1669390400
transform 1 0 8512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_77
timestamp 1669390400
transform 1 0 9968 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_90
timestamp 1669390400
transform 1 0 11424 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_94
timestamp 1669390400
transform 1 0 11872 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_115
timestamp 1669390400
transform 1 0 14224 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_117
timestamp 1669390400
transform 1 0 14448 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_124
timestamp 1669390400
transform 1 0 15232 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_134
timestamp 1669390400
transform 1 0 16352 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_138
timestamp 1669390400
transform 1 0 16800 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_147
timestamp 1669390400
transform 1 0 17808 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_151
timestamp 1669390400
transform 1 0 18256 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_158
timestamp 1669390400
transform 1 0 19040 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_167
timestamp 1669390400
transform 1 0 20048 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_189
timestamp 1669390400
transform 1 0 22512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_193
timestamp 1669390400
transform 1 0 22960 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_195
timestamp 1669390400
transform 1 0 23184 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_205
timestamp 1669390400
transform 1 0 24304 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_212
timestamp 1669390400
transform 1 0 25088 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_221
timestamp 1669390400
transform 1 0 26096 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_228
timestamp 1669390400
transform 1 0 26880 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_235
timestamp 1669390400
transform 1 0 27664 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_239
timestamp 1669390400
transform 1 0 28112 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_246
timestamp 1669390400
transform 1 0 28896 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_256
timestamp 1669390400
transform 1 0 30016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_263
timestamp 1669390400
transform 1 0 30800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_267
timestamp 1669390400
transform 1 0 31248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_269
timestamp 1669390400
transform 1 0 31472 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_275
timestamp 1669390400
transform 1 0 32144 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_282
timestamp 1669390400
transform 1 0 32928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_286
timestamp 1669390400
transform 1 0 33376 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_288
timestamp 1669390400
transform 1 0 33600 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_330
timestamp 1669390400
transform 1 0 38304 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_340
timestamp 1669390400
transform 1 0 39424 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_344
timestamp 1669390400
transform 1 0 39872 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_350
timestamp 1669390400
transform 1 0 40544 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_354
timestamp 1669390400
transform 1 0 40992 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_358
timestamp 1669390400
transform 1 0 41440 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_362
timestamp 1669390400
transform 1 0 41888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_7
timestamp 1669390400
transform 1 0 2128 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_15
timestamp 1669390400
transform 1 0 3024 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_25
timestamp 1669390400
transform 1 0 4144 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_31
timestamp 1669390400
transform 1 0 4816 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_40
timestamp 1669390400
transform 1 0 5824 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_42
timestamp 1669390400
transform 1 0 6048 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_45
timestamp 1669390400
transform 1 0 6384 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_55
timestamp 1669390400
transform 1 0 7504 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_57
timestamp 1669390400
transform 1 0 7728 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_65
timestamp 1669390400
transform 1 0 8624 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_67
timestamp 1669390400
transform 1 0 8848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_82
timestamp 1669390400
transform 1 0 10528 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_88
timestamp 1669390400
transform 1 0 11200 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_140
timestamp 1669390400
transform 1 0 17024 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_150
timestamp 1669390400
transform 1 0 18144 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_157
timestamp 1669390400
transform 1 0 18928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_190
timestamp 1669390400
transform 1 0 22624 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_201
timestamp 1669390400
transform 1 0 23856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_211
timestamp 1669390400
transform 1 0 24976 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_221
timestamp 1669390400
transform 1 0 26096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_254
timestamp 1669390400
transform 1 0 29792 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_260
timestamp 1669390400
transform 1 0 30464 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_266
timestamp 1669390400
transform 1 0 31136 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_272
timestamp 1669390400
transform 1 0 31808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_276
timestamp 1669390400
transform 1 0 32256 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_289
timestamp 1669390400
transform 1 0 33712 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_293
timestamp 1669390400
transform 1 0 34160 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_297
timestamp 1669390400
transform 1 0 34608 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_301
timestamp 1669390400
transform 1 0 35056 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_303
timestamp 1669390400
transform 1 0 35280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_308
timestamp 1669390400
transform 1 0 35840 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_312
timestamp 1669390400
transform 1 0 36288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_316
timestamp 1669390400
transform 1 0 36736 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_320
timestamp 1669390400
transform 1 0 37184 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_324
timestamp 1669390400
transform 1 0 37632 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_329
timestamp 1669390400
transform 1 0 38192 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_333
timestamp 1669390400
transform 1 0 38640 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_337
timestamp 1669390400
transform 1 0 39088 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_343
timestamp 1669390400
transform 1 0 39760 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_347
timestamp 1669390400
transform 1 0 40208 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_351
timestamp 1669390400
transform 1 0 40656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_360
timestamp 1669390400
transform 1 0 41664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_362
timestamp 1669390400
transform 1 0 41888 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_365
timestamp 1669390400
transform 1 0 42224 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_10
timestamp 1669390400
transform 1 0 2464 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_18
timestamp 1669390400
transform 1 0 3360 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_26
timestamp 1669390400
transform 1 0 4256 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_44
timestamp 1669390400
transform 1 0 6272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_48
timestamp 1669390400
transform 1 0 6720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_58
timestamp 1669390400
transform 1 0 7840 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_68
timestamp 1669390400
transform 1 0 8960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_72
timestamp 1669390400
transform 1 0 9408 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_102
timestamp 1669390400
transform 1 0 12768 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_112
timestamp 1669390400
transform 1 0 13888 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1669390400
transform 1 0 15232 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_134
timestamp 1669390400
transform 1 0 16352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_143
timestamp 1669390400
transform 1 0 17360 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_151
timestamp 1669390400
transform 1 0 18256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_155
timestamp 1669390400
transform 1 0 18704 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_161
timestamp 1669390400
transform 1 0 19376 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_171
timestamp 1669390400
transform 1 0 20496 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_173
timestamp 1669390400
transform 1 0 20720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_185
timestamp 1669390400
transform 1 0 22064 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_192
timestamp 1669390400
transform 1 0 22848 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_194
timestamp 1669390400
transform 1 0 23072 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_202
timestamp 1669390400
transform 1 0 23968 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_204
timestamp 1669390400
transform 1 0 24192 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_213
timestamp 1669390400
transform 1 0 25200 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_219
timestamp 1669390400
transform 1 0 25872 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_229
timestamp 1669390400
transform 1 0 26992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_236
timestamp 1669390400
transform 1 0 27776 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_255
timestamp 1669390400
transform 1 0 29904 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_261
timestamp 1669390400
transform 1 0 30576 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_267
timestamp 1669390400
transform 1 0 31248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_273
timestamp 1669390400
transform 1 0 31920 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_279
timestamp 1669390400
transform 1 0 32592 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_283
timestamp 1669390400
transform 1 0 33040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_287
timestamp 1669390400
transform 1 0 33488 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_291
timestamp 1669390400
transform 1 0 33936 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_295
timestamp 1669390400
transform 1 0 34384 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_299
timestamp 1669390400
transform 1 0 34832 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_303
timestamp 1669390400
transform 1 0 35280 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_307
timestamp 1669390400
transform 1 0 35728 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_311
timestamp 1669390400
transform 1 0 36176 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_315
timestamp 1669390400
transform 1 0 36624 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_324
timestamp 1669390400
transform 1 0 37632 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_328 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38080 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_360
timestamp 1669390400
transform 1 0 41664 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_364
timestamp 1669390400
transform 1 0 42112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_33
timestamp 1669390400
transform 1 0 5040 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_41
timestamp 1669390400
transform 1 0 5936 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_48
timestamp 1669390400
transform 1 0 6720 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_56
timestamp 1669390400
transform 1 0 7616 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_63
timestamp 1669390400
transform 1 0 8400 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_84
timestamp 1669390400
transform 1 0 10752 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_86
timestamp 1669390400
transform 1 0 10976 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_89
timestamp 1669390400
transform 1 0 11312 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_96
timestamp 1669390400
transform 1 0 12096 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_103
timestamp 1669390400
transform 1 0 12880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_110
timestamp 1669390400
transform 1 0 13664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_114
timestamp 1669390400
transform 1 0 14112 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_122
timestamp 1669390400
transform 1 0 15008 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_131
timestamp 1669390400
transform 1 0 16016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_135
timestamp 1669390400
transform 1 0 16464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_146
timestamp 1669390400
transform 1 0 17696 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_152
timestamp 1669390400
transform 1 0 18368 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_159
timestamp 1669390400
transform 1 0 19152 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_166
timestamp 1669390400
transform 1 0 19936 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_173
timestamp 1669390400
transform 1 0 20720 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_177
timestamp 1669390400
transform 1 0 21168 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_187
timestamp 1669390400
transform 1 0 22288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_193
timestamp 1669390400
transform 1 0 22960 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_203
timestamp 1669390400
transform 1 0 24080 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_210
timestamp 1669390400
transform 1 0 24864 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_218
timestamp 1669390400
transform 1 0 25760 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_228
timestamp 1669390400
transform 1 0 26880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_235
timestamp 1669390400
transform 1 0 27664 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_242
timestamp 1669390400
transform 1 0 28448 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_248
timestamp 1669390400
transform 1 0 29120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_252
timestamp 1669390400
transform 1 0 29568 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_256
timestamp 1669390400
transform 1 0 30016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_260
timestamp 1669390400
transform 1 0 30464 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_264
timestamp 1669390400
transform 1 0 30912 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_268
timestamp 1669390400
transform 1 0 31360 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_272
timestamp 1669390400
transform 1 0 31808 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_274
timestamp 1669390400
transform 1 0 32032 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_277
timestamp 1669390400
transform 1 0 32368 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_281
timestamp 1669390400
transform 1 0 32816 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_289
timestamp 1669390400
transform 1 0 33712 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_293
timestamp 1669390400
transform 1 0 34160 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_297
timestamp 1669390400
transform 1 0 34608 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_301
timestamp 1669390400
transform 1 0 35056 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_305
timestamp 1669390400
transform 1 0 35504 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_309
timestamp 1669390400
transform 1 0 35952 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_341 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 39536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_349
timestamp 1669390400
transform 1 0 40432 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1669390400
transform 1 0 40880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_365
timestamp 1669390400
transform 1 0 42224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_12
timestamp 1669390400
transform 1 0 2688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_16
timestamp 1669390400
transform 1 0 3136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_23
timestamp 1669390400
transform 1 0 3920 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1669390400
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_44
timestamp 1669390400
transform 1 0 6272 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_46
timestamp 1669390400
transform 1 0 6496 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_49
timestamp 1669390400
transform 1 0 6832 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_56
timestamp 1669390400
transform 1 0 7616 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_63
timestamp 1669390400
transform 1 0 8400 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_94
timestamp 1669390400
transform 1 0 11872 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_98
timestamp 1669390400
transform 1 0 12320 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_117
timestamp 1669390400
transform 1 0 14448 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_127
timestamp 1669390400
transform 1 0 15568 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_135
timestamp 1669390400
transform 1 0 16464 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_144
timestamp 1669390400
transform 1 0 17472 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_154
timestamp 1669390400
transform 1 0 18592 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_158
timestamp 1669390400
transform 1 0 19040 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_164
timestamp 1669390400
transform 1 0 19712 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_173
timestamp 1669390400
transform 1 0 20720 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_188
timestamp 1669390400
transform 1 0 22400 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_221
timestamp 1669390400
transform 1 0 26096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_230
timestamp 1669390400
transform 1 0 27104 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_236
timestamp 1669390400
transform 1 0 27776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_240
timestamp 1669390400
transform 1 0 28224 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_244
timestamp 1669390400
transform 1 0 28672 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_253
timestamp 1669390400
transform 1 0 29680 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_257
timestamp 1669390400
transform 1 0 30128 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_261
timestamp 1669390400
transform 1 0 30576 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_265
timestamp 1669390400
transform 1 0 31024 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_271
timestamp 1669390400
transform 1 0 31696 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_275
timestamp 1669390400
transform 1 0 32144 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_279
timestamp 1669390400
transform 1 0 32592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_283
timestamp 1669390400
transform 1 0 33040 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_287
timestamp 1669390400
transform 1 0 33488 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_291
timestamp 1669390400
transform 1 0 33936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_293
timestamp 1669390400
transform 1 0 34160 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_296 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 34496 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_312
timestamp 1669390400
transform 1 0 36288 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_316
timestamp 1669390400
transform 1 0 36736 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_353
timestamp 1669390400
transform 1 0 40880 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_361
timestamp 1669390400
transform 1 0 41776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_365
timestamp 1669390400
transform 1 0 42224 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_9
timestamp 1669390400
transform 1 0 2352 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_16
timestamp 1669390400
transform 1 0 3136 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_23
timestamp 1669390400
transform 1 0 3920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_30
timestamp 1669390400
transform 1 0 4704 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_37
timestamp 1669390400
transform 1 0 5488 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_47
timestamp 1669390400
transform 1 0 6608 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_49
timestamp 1669390400
transform 1 0 6832 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_57
timestamp 1669390400
transform 1 0 7728 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_68
timestamp 1669390400
transform 1 0 8960 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_75
timestamp 1669390400
transform 1 0 9744 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_81
timestamp 1669390400
transform 1 0 10416 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_88
timestamp 1669390400
transform 1 0 11200 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_95
timestamp 1669390400
transform 1 0 11984 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_104
timestamp 1669390400
transform 1 0 12992 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_112
timestamp 1669390400
transform 1 0 13888 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_116
timestamp 1669390400
transform 1 0 14336 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_126
timestamp 1669390400
transform 1 0 15456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_136
timestamp 1669390400
transform 1 0 16576 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_138
timestamp 1669390400
transform 1 0 16800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_150
timestamp 1669390400
transform 1 0 18144 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_160
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_166
timestamp 1669390400
transform 1 0 19936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_175
timestamp 1669390400
transform 1 0 20944 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_184
timestamp 1669390400
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_196
timestamp 1669390400
transform 1 0 23296 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_202
timestamp 1669390400
transform 1 0 23968 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_209
timestamp 1669390400
transform 1 0 24752 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_220
timestamp 1669390400
transform 1 0 25984 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_224
timestamp 1669390400
transform 1 0 26432 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_228
timestamp 1669390400
transform 1 0 26880 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_232
timestamp 1669390400
transform 1 0 27328 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_236
timestamp 1669390400
transform 1 0 27776 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_240
timestamp 1669390400
transform 1 0 28224 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_244
timestamp 1669390400
transform 1 0 28672 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_248
timestamp 1669390400
transform 1 0 29120 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_252
timestamp 1669390400
transform 1 0 29568 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_256
timestamp 1669390400
transform 1 0 30016 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_260
timestamp 1669390400
transform 1 0 30464 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_264
timestamp 1669390400
transform 1 0 30912 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_268
timestamp 1669390400
transform 1 0 31360 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_272
timestamp 1669390400
transform 1 0 31808 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_276
timestamp 1669390400
transform 1 0 32256 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_280
timestamp 1669390400
transform 1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_365
timestamp 1669390400
transform 1 0 42224 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_5
timestamp 1669390400
transform 1 0 1904 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_12
timestamp 1669390400
transform 1 0 2688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_19
timestamp 1669390400
transform 1 0 3472 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_26
timestamp 1669390400
transform 1 0 4256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_44
timestamp 1669390400
transform 1 0 6272 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_53
timestamp 1669390400
transform 1 0 7280 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_84
timestamp 1669390400
transform 1 0 10752 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_91
timestamp 1669390400
transform 1 0 11536 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_98
timestamp 1669390400
transform 1 0 12320 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_115
timestamp 1669390400
transform 1 0 14224 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_122
timestamp 1669390400
transform 1 0 15008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_130
timestamp 1669390400
transform 1 0 15904 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_137
timestamp 1669390400
transform 1 0 16688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_145
timestamp 1669390400
transform 1 0 17584 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_152
timestamp 1669390400
transform 1 0 18368 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_158
timestamp 1669390400
transform 1 0 19040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_165
timestamp 1669390400
transform 1 0 19824 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_174
timestamp 1669390400
transform 1 0 20832 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_187
timestamp 1669390400
transform 1 0 22288 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_193
timestamp 1669390400
transform 1 0 22960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_197
timestamp 1669390400
transform 1 0 23408 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_201
timestamp 1669390400
transform 1 0 23856 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_204
timestamp 1669390400
transform 1 0 24192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_208
timestamp 1669390400
transform 1 0 24640 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_211
timestamp 1669390400
transform 1 0 24976 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_215
timestamp 1669390400
transform 1 0 25424 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_221
timestamp 1669390400
transform 1 0 26096 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_225
timestamp 1669390400
transform 1 0 26544 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_229
timestamp 1669390400
transform 1 0 26992 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_233
timestamp 1669390400
transform 1 0 27440 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_237
timestamp 1669390400
transform 1 0 27888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_241
timestamp 1669390400
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_253
timestamp 1669390400
transform 1 0 29680 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_257
timestamp 1669390400
transform 1 0 30128 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_289
timestamp 1669390400
transform 1 0 33712 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_305
timestamp 1669390400
transform 1 0 35504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_313
timestamp 1669390400
transform 1 0 36400 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_317
timestamp 1669390400
transform 1 0 36848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_353
timestamp 1669390400
transform 1 0 40880 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_361
timestamp 1669390400
transform 1 0 41776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_365
timestamp 1669390400
transform 1 0 42224 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_9
timestamp 1669390400
transform 1 0 2352 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_16
timestamp 1669390400
transform 1 0 3136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_24
timestamp 1669390400
transform 1 0 4032 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_31
timestamp 1669390400
transform 1 0 4816 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_38
timestamp 1669390400
transform 1 0 5600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_42
timestamp 1669390400
transform 1 0 6048 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_48
timestamp 1669390400
transform 1 0 6720 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_52
timestamp 1669390400
transform 1 0 7168 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_59
timestamp 1669390400
transform 1 0 7952 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_76
timestamp 1669390400
transform 1 0 9856 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_83
timestamp 1669390400
transform 1 0 10640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_87
timestamp 1669390400
transform 1 0 11088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_97
timestamp 1669390400
transform 1 0 12208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_104
timestamp 1669390400
transform 1 0 12992 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_116
timestamp 1669390400
transform 1 0 14336 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_126
timestamp 1669390400
transform 1 0 15456 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_128
timestamp 1669390400
transform 1 0 15680 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_131
timestamp 1669390400
transform 1 0 16016 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_138
timestamp 1669390400
transform 1 0 16800 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_149
timestamp 1669390400
transform 1 0 18032 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_156
timestamp 1669390400
transform 1 0 18816 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_160
timestamp 1669390400
transform 1 0 19264 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_162
timestamp 1669390400
transform 1 0 19488 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_168
timestamp 1669390400
transform 1 0 20160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_172
timestamp 1669390400
transform 1 0 20608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_175
timestamp 1669390400
transform 1 0 20944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_177
timestamp 1669390400
transform 1 0 21168 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_180
timestamp 1669390400
transform 1 0 21504 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_184
timestamp 1669390400
transform 1 0 21952 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_188
timestamp 1669390400
transform 1 0 22400 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_192
timestamp 1669390400
transform 1 0 22848 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_196
timestamp 1669390400
transform 1 0 23296 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_200
timestamp 1669390400
transform 1 0 23744 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_204
timestamp 1669390400
transform 1 0 24192 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_207
timestamp 1669390400
transform 1 0 24528 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_211
timestamp 1669390400
transform 1 0 24976 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_218
timestamp 1669390400
transform 1 0 25760 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_222
timestamp 1669390400
transform 1 0 26208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_226
timestamp 1669390400
transform 1 0 26656 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_230
timestamp 1669390400
transform 1 0 27104 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_234
timestamp 1669390400
transform 1 0 27552 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_238
timestamp 1669390400
transform 1 0 28000 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_270
timestamp 1669390400
transform 1 0 31584 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_278
timestamp 1669390400
transform 1 0 32480 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_282
timestamp 1669390400
transform 1 0 32928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_365
timestamp 1669390400
transform 1 0 42224 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_8
timestamp 1669390400
transform 1 0 2240 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_12
timestamp 1669390400
transform 1 0 2688 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_16
timestamp 1669390400
transform 1 0 3136 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_20
timestamp 1669390400
transform 1 0 3584 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_26
timestamp 1669390400
transform 1 0 4256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_28
timestamp 1669390400
transform 1 0 4480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_40
timestamp 1669390400
transform 1 0 5824 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_47
timestamp 1669390400
transform 1 0 6608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_51
timestamp 1669390400
transform 1 0 7056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_57
timestamp 1669390400
transform 1 0 7728 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_66
timestamp 1669390400
transform 1 0 8736 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_97
timestamp 1669390400
transform 1 0 12208 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_110
timestamp 1669390400
transform 1 0 13664 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_116
timestamp 1669390400
transform 1 0 14336 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_123
timestamp 1669390400
transform 1 0 15120 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_127
timestamp 1669390400
transform 1 0 15568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_133
timestamp 1669390400
transform 1 0 16240 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_137
timestamp 1669390400
transform 1 0 16688 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_140
timestamp 1669390400
transform 1 0 17024 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_142
timestamp 1669390400
transform 1 0 17248 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_145
timestamp 1669390400
transform 1 0 17584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_151
timestamp 1669390400
transform 1 0 18256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_155
timestamp 1669390400
transform 1 0 18704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_159
timestamp 1669390400
transform 1 0 19152 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_163
timestamp 1669390400
transform 1 0 19600 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_165
timestamp 1669390400
transform 1 0 19824 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_168
timestamp 1669390400
transform 1 0 20160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_182
timestamp 1669390400
transform 1 0 21728 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_186
timestamp 1669390400
transform 1 0 22176 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_188
timestamp 1669390400
transform 1 0 22400 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_191
timestamp 1669390400
transform 1 0 22736 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_195
timestamp 1669390400
transform 1 0 23184 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_197
timestamp 1669390400
transform 1 0 23408 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_200
timestamp 1669390400
transform 1 0 23744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_204
timestamp 1669390400
transform 1 0 24192 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_207
timestamp 1669390400
transform 1 0 24528 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_223
timestamp 1669390400
transform 1 0 26320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_229
timestamp 1669390400
transform 1 0 26992 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_245
timestamp 1669390400
transform 1 0 28784 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_353
timestamp 1669390400
transform 1 0 40880 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_361
timestamp 1669390400
transform 1 0 41776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_365
timestamp 1669390400
transform 1 0 42224 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_5
timestamp 1669390400
transform 1 0 1904 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_9
timestamp 1669390400
transform 1 0 2352 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_13
timestamp 1669390400
transform 1 0 2800 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_17
timestamp 1669390400
transform 1 0 3248 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_21
timestamp 1669390400
transform 1 0 3696 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_25
timestamp 1669390400
transform 1 0 4144 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_29
timestamp 1669390400
transform 1 0 4592 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_33
timestamp 1669390400
transform 1 0 5040 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_37
timestamp 1669390400
transform 1 0 5488 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_41
timestamp 1669390400
transform 1 0 5936 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_48
timestamp 1669390400
transform 1 0 6720 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_50
timestamp 1669390400
transform 1 0 6944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_56
timestamp 1669390400
transform 1 0 7616 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_63
timestamp 1669390400
transform 1 0 8400 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_79
timestamp 1669390400
transform 1 0 10192 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_88
timestamp 1669390400
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_94
timestamp 1669390400
transform 1 0 11872 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_98
timestamp 1669390400
transform 1 0 12320 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_105
timestamp 1669390400
transform 1 0 13104 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_111
timestamp 1669390400
transform 1 0 13776 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_117
timestamp 1669390400
transform 1 0 14448 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_121
timestamp 1669390400
transform 1 0 14896 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_125
timestamp 1669390400
transform 1 0 15344 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_129
timestamp 1669390400
transform 1 0 15792 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_131
timestamp 1669390400
transform 1 0 16016 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_134
timestamp 1669390400
transform 1 0 16352 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_138
timestamp 1669390400
transform 1 0 16800 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_147
timestamp 1669390400
transform 1 0 17808 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_149
timestamp 1669390400
transform 1 0 18032 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_152
timestamp 1669390400
transform 1 0 18368 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_156
timestamp 1669390400
transform 1 0 18816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_160
timestamp 1669390400
transform 1 0 19264 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_162
timestamp 1669390400
transform 1 0 19488 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_165
timestamp 1669390400
transform 1 0 19824 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1669390400
transform 1 0 20272 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_173
timestamp 1669390400
transform 1 0 20720 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_177
timestamp 1669390400
transform 1 0 21168 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_179
timestamp 1669390400
transform 1 0 21392 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_182
timestamp 1669390400
transform 1 0 21728 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_186
timestamp 1669390400
transform 1 0 22176 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_190
timestamp 1669390400
transform 1 0 22624 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_194
timestamp 1669390400
transform 1 0 23072 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_210
timestamp 1669390400
transform 1 0 24864 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_365
timestamp 1669390400
transform 1 0 42224 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_6
timestamp 1669390400
transform 1 0 2016 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_10
timestamp 1669390400
transform 1 0 2464 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_14
timestamp 1669390400
transform 1 0 2912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_18
timestamp 1669390400
transform 1 0 3360 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_22
timestamp 1669390400
transform 1 0 3808 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_26
timestamp 1669390400
transform 1 0 4256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_30
timestamp 1669390400
transform 1 0 4704 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_41
timestamp 1669390400
transform 1 0 5936 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_45
timestamp 1669390400
transform 1 0 6384 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_49
timestamp 1669390400
transform 1 0 6832 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_53
timestamp 1669390400
transform 1 0 7280 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_57
timestamp 1669390400
transform 1 0 7728 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_63
timestamp 1669390400
transform 1 0 8400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_65
timestamp 1669390400
transform 1 0 8624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_70
timestamp 1669390400
transform 1 0 9184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1669390400
transform 1 0 10192 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_83
timestamp 1669390400
transform 1 0 10640 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_87
timestamp 1669390400
transform 1 0 11088 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_90
timestamp 1669390400
transform 1 0 11424 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_94
timestamp 1669390400
transform 1 0 11872 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_96
timestamp 1669390400
transform 1 0 12096 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_99
timestamp 1669390400
transform 1 0 12432 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_103
timestamp 1669390400
transform 1 0 12880 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_111
timestamp 1669390400
transform 1 0 13776 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_113
timestamp 1669390400
transform 1 0 14000 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_116
timestamp 1669390400
transform 1 0 14336 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_120
timestamp 1669390400
transform 1 0 14784 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_124
timestamp 1669390400
transform 1 0 15232 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_128
timestamp 1669390400
transform 1 0 15680 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_132
timestamp 1669390400
transform 1 0 16128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_134
timestamp 1669390400
transform 1 0 16352 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_137
timestamp 1669390400
transform 1 0 16688 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_141
timestamp 1669390400
transform 1 0 17136 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_145
timestamp 1669390400
transform 1 0 17584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_151
timestamp 1669390400
transform 1 0 18256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_155
timestamp 1669390400
transform 1 0 18704 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_159
timestamp 1669390400
transform 1 0 19152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_163
timestamp 1669390400
transform 1 0 19600 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_167
timestamp 1669390400
transform 1 0 20048 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_171
timestamp 1669390400
transform 1 0 20496 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_175
timestamp 1669390400
transform 1 0 20944 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_182
timestamp 1669390400
transform 1 0 21728 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_186
timestamp 1669390400
transform 1 0 22176 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_190
timestamp 1669390400
transform 1 0 22624 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_222
timestamp 1669390400
transform 1 0 26208 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_238
timestamp 1669390400
transform 1 0 28000 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1669390400
transform 1 0 28896 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_353
timestamp 1669390400
transform 1 0 40880 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_361
timestamp 1669390400
transform 1 0 41776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_365
timestamp 1669390400
transform 1 0 42224 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_6
timestamp 1669390400
transform 1 0 2016 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_10
timestamp 1669390400
transform 1 0 2464 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_14
timestamp 1669390400
transform 1 0 2912 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_18
timestamp 1669390400
transform 1 0 3360 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_22
timestamp 1669390400
transform 1 0 3808 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_25
timestamp 1669390400
transform 1 0 4144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_29
timestamp 1669390400
transform 1 0 4592 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_32
timestamp 1669390400
transform 1 0 4928 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_36
timestamp 1669390400
transform 1 0 5376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_40
timestamp 1669390400
transform 1 0 5824 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_43
timestamp 1669390400
transform 1 0 6160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_47
timestamp 1669390400
transform 1 0 6608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_50
timestamp 1669390400
transform 1 0 6944 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_54
timestamp 1669390400
transform 1 0 7392 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_58
timestamp 1669390400
transform 1 0 7840 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_62
timestamp 1669390400
transform 1 0 8288 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_76
timestamp 1669390400
transform 1 0 9856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_80
timestamp 1669390400
transform 1 0 10304 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_83
timestamp 1669390400
transform 1 0 10640 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_87
timestamp 1669390400
transform 1 0 11088 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_91
timestamp 1669390400
transform 1 0 11536 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_97
timestamp 1669390400
transform 1 0 12208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_101
timestamp 1669390400
transform 1 0 12656 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_105
timestamp 1669390400
transform 1 0 13104 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_109
timestamp 1669390400
transform 1 0 13552 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_115
timestamp 1669390400
transform 1 0 14224 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_119
timestamp 1669390400
transform 1 0 14672 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_121
timestamp 1669390400
transform 1 0 14896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_124
timestamp 1669390400
transform 1 0 15232 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_126
timestamp 1669390400
transform 1 0 15456 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_129
timestamp 1669390400
transform 1 0 15792 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_133
timestamp 1669390400
transform 1 0 16240 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_135
timestamp 1669390400
transform 1 0 16464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_138
timestamp 1669390400
transform 1 0 16800 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_146
timestamp 1669390400
transform 1 0 17696 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_149
timestamp 1669390400
transform 1 0 18032 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_153
timestamp 1669390400
transform 1 0 18480 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_157
timestamp 1669390400
transform 1 0 18928 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_161
timestamp 1669390400
transform 1 0 19376 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_165
timestamp 1669390400
transform 1 0 19824 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_169
timestamp 1669390400
transform 1 0 20272 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_173
timestamp 1669390400
transform 1 0 20720 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_177
timestamp 1669390400
transform 1 0 21168 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_181
timestamp 1669390400
transform 1 0 21616 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_365
timestamp 1669390400
transform 1 0 42224 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_4
timestamp 1669390400
transform 1 0 1792 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_7
timestamp 1669390400
transform 1 0 2128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_11
timestamp 1669390400
transform 1 0 2576 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_15
timestamp 1669390400
transform 1 0 3024 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_21
timestamp 1669390400
transform 1 0 3696 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_25
timestamp 1669390400
transform 1 0 4144 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_27
timestamp 1669390400
transform 1 0 4368 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_30
timestamp 1669390400
transform 1 0 4704 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_40
timestamp 1669390400
transform 1 0 5824 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_42
timestamp 1669390400
transform 1 0 6048 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_45
timestamp 1669390400
transform 1 0 6384 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_49
timestamp 1669390400
transform 1 0 6832 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_53
timestamp 1669390400
transform 1 0 7280 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_57
timestamp 1669390400
transform 1 0 7728 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_61
timestamp 1669390400
transform 1 0 8176 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_63
timestamp 1669390400
transform 1 0 8400 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_66
timestamp 1669390400
transform 1 0 8736 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_70
timestamp 1669390400
transform 1 0 9184 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_74
timestamp 1669390400
transform 1 0 9632 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_78
timestamp 1669390400
transform 1 0 10080 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_81
timestamp 1669390400
transform 1 0 10416 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_85
timestamp 1669390400
transform 1 0 10864 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_91
timestamp 1669390400
transform 1 0 11536 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_93
timestamp 1669390400
transform 1 0 11760 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_96
timestamp 1669390400
transform 1 0 12096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_100
timestamp 1669390400
transform 1 0 12544 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_102
timestamp 1669390400
transform 1 0 12768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_111
timestamp 1669390400
transform 1 0 13776 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_113
timestamp 1669390400
transform 1 0 14000 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_116
timestamp 1669390400
transform 1 0 14336 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_120
timestamp 1669390400
transform 1 0 14784 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_124
timestamp 1669390400
transform 1 0 15232 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_130
timestamp 1669390400
transform 1 0 15904 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_134
timestamp 1669390400
transform 1 0 16352 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_138
timestamp 1669390400
transform 1 0 16800 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_142
timestamp 1669390400
transform 1 0 17248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_145
timestamp 1669390400
transform 1 0 17584 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_149
timestamp 1669390400
transform 1 0 18032 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_153
timestamp 1669390400
transform 1 0 18480 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_157
timestamp 1669390400
transform 1 0 18928 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_161
timestamp 1669390400
transform 1 0 19376 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_165
timestamp 1669390400
transform 1 0 19824 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_169
timestamp 1669390400
transform 1 0 20272 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_353
timestamp 1669390400
transform 1 0 40880 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_361
timestamp 1669390400
transform 1 0 41776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_365
timestamp 1669390400
transform 1 0 42224 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_8
timestamp 1669390400
transform 1 0 2240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_12
timestamp 1669390400
transform 1 0 2688 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_16
timestamp 1669390400
transform 1 0 3136 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_20
timestamp 1669390400
transform 1 0 3584 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_24
timestamp 1669390400
transform 1 0 4032 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_28
timestamp 1669390400
transform 1 0 4480 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_32
timestamp 1669390400
transform 1 0 4928 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_34
timestamp 1669390400
transform 1 0 5152 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_37
timestamp 1669390400
transform 1 0 5488 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_41
timestamp 1669390400
transform 1 0 5936 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_45
timestamp 1669390400
transform 1 0 6384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_49
timestamp 1669390400
transform 1 0 6832 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_53
timestamp 1669390400
transform 1 0 7280 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_57
timestamp 1669390400
transform 1 0 7728 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_61
timestamp 1669390400
transform 1 0 8176 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_65
timestamp 1669390400
transform 1 0 8624 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_67
timestamp 1669390400
transform 1 0 8848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_76
timestamp 1669390400
transform 1 0 9856 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_80
timestamp 1669390400
transform 1 0 10304 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_84
timestamp 1669390400
transform 1 0 10752 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_88
timestamp 1669390400
transform 1 0 11200 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_92
timestamp 1669390400
transform 1 0 11648 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_96
timestamp 1669390400
transform 1 0 12096 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_100
timestamp 1669390400
transform 1 0 12544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_104
timestamp 1669390400
transform 1 0 12992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_107
timestamp 1669390400
transform 1 0 13328 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_111
timestamp 1669390400
transform 1 0 13776 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_115
timestamp 1669390400
transform 1 0 14224 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_119
timestamp 1669390400
transform 1 0 14672 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_123
timestamp 1669390400
transform 1 0 15120 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_125
timestamp 1669390400
transform 1 0 15344 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_128
timestamp 1669390400
transform 1 0 15680 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_130
timestamp 1669390400
transform 1 0 15904 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_133
timestamp 1669390400
transform 1 0 16240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_147
timestamp 1669390400
transform 1 0 17808 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_151
timestamp 1669390400
transform 1 0 18256 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_155
timestamp 1669390400
transform 1 0 18704 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_159
timestamp 1669390400
transform 1 0 19152 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_163
timestamp 1669390400
transform 1 0 19600 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_195
timestamp 1669390400
transform 1 0 23184 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_211
timestamp 1669390400
transform 1 0 24976 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_365
timestamp 1669390400
transform 1 0 42224 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_5
timestamp 1669390400
transform 1 0 1904 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_9
timestamp 1669390400
transform 1 0 2352 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_13
timestamp 1669390400
transform 1 0 2800 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_17
timestamp 1669390400
transform 1 0 3248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_21
timestamp 1669390400
transform 1 0 3696 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_25
timestamp 1669390400
transform 1 0 4144 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_29
timestamp 1669390400
transform 1 0 4592 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_33
timestamp 1669390400
transform 1 0 5040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_43
timestamp 1669390400
transform 1 0 6160 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_47
timestamp 1669390400
transform 1 0 6608 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_51
timestamp 1669390400
transform 1 0 7056 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_55
timestamp 1669390400
transform 1 0 7504 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_58
timestamp 1669390400
transform 1 0 7840 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_62
timestamp 1669390400
transform 1 0 8288 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_66
timestamp 1669390400
transform 1 0 8736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_70
timestamp 1669390400
transform 1 0 9184 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_74
timestamp 1669390400
transform 1 0 9632 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_76
timestamp 1669390400
transform 1 0 9856 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_79
timestamp 1669390400
transform 1 0 10192 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_83
timestamp 1669390400
transform 1 0 10640 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_87
timestamp 1669390400
transform 1 0 11088 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_91
timestamp 1669390400
transform 1 0 11536 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_95
timestamp 1669390400
transform 1 0 11984 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_97
timestamp 1669390400
transform 1 0 12208 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_100
timestamp 1669390400
transform 1 0 12544 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_104
timestamp 1669390400
transform 1 0 12992 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_111
timestamp 1669390400
transform 1 0 13776 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_115
timestamp 1669390400
transform 1 0 14224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_119
timestamp 1669390400
transform 1 0 14672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_122
timestamp 1669390400
transform 1 0 15008 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_126
timestamp 1669390400
transform 1 0 15456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_130
timestamp 1669390400
transform 1 0 15904 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_133
timestamp 1669390400
transform 1 0 16240 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_137
timestamp 1669390400
transform 1 0 16688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_141
timestamp 1669390400
transform 1 0 17136 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_145
timestamp 1669390400
transform 1 0 17584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_149
timestamp 1669390400
transform 1 0 18032 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_153
timestamp 1669390400
transform 1 0 18480 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_169
timestamp 1669390400
transform 1 0 20272 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_329
timestamp 1669390400
transform 1 0 38192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_333
timestamp 1669390400
transform 1 0 38640 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_348
timestamp 1669390400
transform 1 0 40320 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_352
timestamp 1669390400
transform 1 0 40768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_360
timestamp 1669390400
transform 1 0 41664 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_364
timestamp 1669390400
transform 1 0 42112 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_5
timestamp 1669390400
transform 1 0 1904 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_9
timestamp 1669390400
transform 1 0 2352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_13
timestamp 1669390400
transform 1 0 2800 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1669390400
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_21
timestamp 1669390400
transform 1 0 3696 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_25
timestamp 1669390400
transform 1 0 4144 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_29
timestamp 1669390400
transform 1 0 4592 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_33
timestamp 1669390400
transform 1 0 5040 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_35
timestamp 1669390400
transform 1 0 5264 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_38
timestamp 1669390400
transform 1 0 5600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_44
timestamp 1669390400
transform 1 0 6272 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_48
timestamp 1669390400
transform 1 0 6720 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_52
timestamp 1669390400
transform 1 0 7168 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_56
timestamp 1669390400
transform 1 0 7616 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_60
timestamp 1669390400
transform 1 0 8064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_76
timestamp 1669390400
transform 1 0 9856 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_80
timestamp 1669390400
transform 1 0 10304 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_84
timestamp 1669390400
transform 1 0 10752 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_90
timestamp 1669390400
transform 1 0 11424 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_96
timestamp 1669390400
transform 1 0 12096 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_100
timestamp 1669390400
transform 1 0 12544 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_102
timestamp 1669390400
transform 1 0 12768 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_105
timestamp 1669390400
transform 1 0 13104 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_109
timestamp 1669390400
transform 1 0 13552 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_113
timestamp 1669390400
transform 1 0 14000 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_117
timestamp 1669390400
transform 1 0 14448 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_120
timestamp 1669390400
transform 1 0 14784 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_124
timestamp 1669390400
transform 1 0 15232 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_128
timestamp 1669390400
transform 1 0 15680 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_132
timestamp 1669390400
transform 1 0 16128 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_136
timestamp 1669390400
transform 1 0 16576 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_140
timestamp 1669390400
transform 1 0 17024 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_365
timestamp 1669390400
transform 1 0 42224 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_6
timestamp 1669390400
transform 1 0 2016 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_10
timestamp 1669390400
transform 1 0 2464 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_14
timestamp 1669390400
transform 1 0 2912 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_18
timestamp 1669390400
transform 1 0 3360 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_22
timestamp 1669390400
transform 1 0 3808 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_26
timestamp 1669390400
transform 1 0 4256 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_30
timestamp 1669390400
transform 1 0 4704 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_40
timestamp 1669390400
transform 1 0 5824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_46
timestamp 1669390400
transform 1 0 6496 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_50
timestamp 1669390400
transform 1 0 6944 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_52
timestamp 1669390400
transform 1 0 7168 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_55
timestamp 1669390400
transform 1 0 7504 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_59
timestamp 1669390400
transform 1 0 7952 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_63
timestamp 1669390400
transform 1 0 8400 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_67
timestamp 1669390400
transform 1 0 8848 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_71
timestamp 1669390400
transform 1 0 9296 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_75
timestamp 1669390400
transform 1 0 9744 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_79
timestamp 1669390400
transform 1 0 10192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_83
timestamp 1669390400
transform 1 0 10640 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_86
timestamp 1669390400
transform 1 0 10976 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_90
timestamp 1669390400
transform 1 0 11424 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_92
timestamp 1669390400
transform 1 0 11648 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_95
timestamp 1669390400
transform 1 0 11984 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_99
timestamp 1669390400
transform 1 0 12432 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_103
timestamp 1669390400
transform 1 0 12880 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_111
timestamp 1669390400
transform 1 0 13776 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_115
timestamp 1669390400
transform 1 0 14224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_119
timestamp 1669390400
transform 1 0 14672 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_123
timestamp 1669390400
transform 1 0 15120 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_155
timestamp 1669390400
transform 1 0 18704 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_171
timestamp 1669390400
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_175
timestamp 1669390400
transform 1 0 20944 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_353
timestamp 1669390400
transform 1 0 40880 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_361
timestamp 1669390400
transform 1 0 41776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_365
timestamp 1669390400
transform 1 0 42224 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_5
timestamp 1669390400
transform 1 0 1904 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_9
timestamp 1669390400
transform 1 0 2352 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_11
timestamp 1669390400
transform 1 0 2576 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_14
timestamp 1669390400
transform 1 0 2912 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_18
timestamp 1669390400
transform 1 0 3360 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_22
timestamp 1669390400
transform 1 0 3808 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_25
timestamp 1669390400
transform 1 0 4144 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_29
timestamp 1669390400
transform 1 0 4592 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_31
timestamp 1669390400
transform 1 0 4816 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_34
timestamp 1669390400
transform 1 0 5152 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_38
timestamp 1669390400
transform 1 0 5600 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_42
timestamp 1669390400
transform 1 0 6048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_46
timestamp 1669390400
transform 1 0 6496 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_50
timestamp 1669390400
transform 1 0 6944 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_54
timestamp 1669390400
transform 1 0 7392 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_58
timestamp 1669390400
transform 1 0 7840 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_62
timestamp 1669390400
transform 1 0 8288 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_75
timestamp 1669390400
transform 1 0 9744 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_78
timestamp 1669390400
transform 1 0 10080 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_82
timestamp 1669390400
transform 1 0 10528 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_85
timestamp 1669390400
transform 1 0 10864 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_89
timestamp 1669390400
transform 1 0 11312 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_121
timestamp 1669390400
transform 1 0 14896 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_365
timestamp 1669390400
transform 1 0 42224 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_6
timestamp 1669390400
transform 1 0 2016 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_8
timestamp 1669390400
transform 1 0 2240 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_11
timestamp 1669390400
transform 1 0 2576 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_15
timestamp 1669390400
transform 1 0 3024 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_31
timestamp 1669390400
transform 1 0 4816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_40
timestamp 1669390400
transform 1 0 5824 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_44
timestamp 1669390400
transform 1 0 6272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_48
timestamp 1669390400
transform 1 0 6720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_51
timestamp 1669390400
transform 1 0 7056 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_55
timestamp 1669390400
transform 1 0 7504 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_59
timestamp 1669390400
transform 1 0 7952 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_67
timestamp 1669390400
transform 1 0 8848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_71
timestamp 1669390400
transform 1 0 9296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_74
timestamp 1669390400
transform 1 0 9632 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_353
timestamp 1669390400
transform 1 0 40880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_361
timestamp 1669390400
transform 1 0 41776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_365
timestamp 1669390400
transform 1 0 42224 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_365
timestamp 1669390400
transform 1 0 42224 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_353
timestamp 1669390400
transform 1 0 40880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_361
timestamp 1669390400
transform 1 0 41776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_365
timestamp 1669390400
transform 1 0 42224 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_365
timestamp 1669390400
transform 1 0 42224 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_353
timestamp 1669390400
transform 1 0 40880 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_361
timestamp 1669390400
transform 1 0 41776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_365
timestamp 1669390400
transform 1 0 42224 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_365
timestamp 1669390400
transform 1 0 42224 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_353
timestamp 1669390400
transform 1 0 40880 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_361
timestamp 1669390400
transform 1 0 41776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_365
timestamp 1669390400
transform 1 0 42224 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_365
timestamp 1669390400
transform 1 0 42224 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_353
timestamp 1669390400
transform 1 0 40880 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_361
timestamp 1669390400
transform 1 0 41776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_365
timestamp 1669390400
transform 1 0 42224 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_365
timestamp 1669390400
transform 1 0 42224 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_353
timestamp 1669390400
transform 1 0 40880 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_361
timestamp 1669390400
transform 1 0 41776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_365
timestamp 1669390400
transform 1 0 42224 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_365
timestamp 1669390400
transform 1 0 42224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_353
timestamp 1669390400
transform 1 0 40880 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_361
timestamp 1669390400
transform 1 0 41776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_365
timestamp 1669390400
transform 1 0 42224 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_365
timestamp 1669390400
transform 1 0 42224 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_353
timestamp 1669390400
transform 1 0 40880 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_361
timestamp 1669390400
transform 1 0 41776 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_365
timestamp 1669390400
transform 1 0 42224 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_365
timestamp 1669390400
transform 1 0 42224 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_353
timestamp 1669390400
transform 1 0 40880 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_361
timestamp 1669390400
transform 1 0 41776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_365
timestamp 1669390400
transform 1 0 42224 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_353
timestamp 1669390400
transform 1 0 40880 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_361
timestamp 1669390400
transform 1 0 41776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_365
timestamp 1669390400
transform 1 0 42224 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_34
timestamp 1669390400
transform 1 0 5152 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_37
timestamp 1669390400
transform 1 0 5488 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_69
timestamp 1669390400
transform 1 0 9072 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_72
timestamp 1669390400
transform 1 0 9408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_104
timestamp 1669390400
transform 1 0 12992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_107
timestamp 1669390400
transform 1 0 13328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_139
timestamp 1669390400
transform 1 0 16912 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_142
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_174
timestamp 1669390400
transform 1 0 20832 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_177
timestamp 1669390400
transform 1 0 21168 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_209
timestamp 1669390400
transform 1 0 24752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_244
timestamp 1669390400
transform 1 0 28672 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_247
timestamp 1669390400
transform 1 0 29008 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_282
timestamp 1669390400
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_314
timestamp 1669390400
transform 1 0 36512 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_317
timestamp 1669390400
transform 1 0 36848 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_349
timestamp 1669390400
transform 1 0 40432 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_352
timestamp 1669390400
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_360
timestamp 1669390400
transform 1 0 41664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_364
timestamp 1669390400
transform 1 0 42112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 42560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 42560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 42560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 42560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 42560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 42560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 42560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 42560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 42560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 42560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 42560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 42560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 42560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 42560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 42560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 42560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 42560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 42560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 42560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 42560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 42560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 42560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 42560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 42560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 42560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 42560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 5264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 13104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 20944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 28784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 36624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _344_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14560 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _345_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13552 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _346_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15792 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _347_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 14560 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _348_
timestamp 1669390400
transform 1 0 40544 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _349_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _350_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _351_
timestamp 1669390400
transform 1 0 5600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _352_
timestamp 1669390400
transform 1 0 10864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _353_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17472 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _354_
timestamp 1669390400
transform 1 0 27328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _355_
timestamp 1669390400
transform -1 0 24752 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _356_
timestamp 1669390400
transform 1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _357_
timestamp 1669390400
transform 1 0 28672 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _358_
timestamp 1669390400
transform -1 0 33040 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _359_
timestamp 1669390400
transform 1 0 10976 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _360_
timestamp 1669390400
transform 1 0 11424 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _361_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26096 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _362_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29008 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _363_
timestamp 1669390400
transform 1 0 31248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _364_
timestamp 1669390400
transform -1 0 34160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _365_
timestamp 1669390400
transform -1 0 31808 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _366_
timestamp 1669390400
transform -1 0 34160 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _367_
timestamp 1669390400
transform -1 0 31920 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1669390400
transform 1 0 31696 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _369_
timestamp 1669390400
transform -1 0 35840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _370_
timestamp 1669390400
transform 1 0 34384 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _371_
timestamp 1669390400
transform 1 0 38080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _372_
timestamp 1669390400
transform -1 0 40432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _373_
timestamp 1669390400
transform 1 0 33264 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1669390400
transform -1 0 42112 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _375_
timestamp 1669390400
transform 1 0 41776 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _376_
timestamp 1669390400
transform -1 0 42112 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _377_
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _378_
timestamp 1669390400
transform 1 0 41440 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _379_
timestamp 1669390400
transform -1 0 40432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _380_
timestamp 1669390400
transform -1 0 39760 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _381_
timestamp 1669390400
transform 1 0 37744 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _382_
timestamp 1669390400
transform 1 0 41440 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _383_
timestamp 1669390400
transform 1 0 39424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _384_
timestamp 1669390400
transform 1 0 39984 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _385_
timestamp 1669390400
transform -1 0 12992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _386_
timestamp 1669390400
transform 1 0 7056 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _387_
timestamp 1669390400
transform -1 0 11872 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _388_
timestamp 1669390400
transform 1 0 6160 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _389_
timestamp 1669390400
transform 1 0 8288 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _390_
timestamp 1669390400
transform -1 0 2688 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _391_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _392_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11200 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _393_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 14896 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _394_
timestamp 1669390400
transform -1 0 10976 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _395_
timestamp 1669390400
transform -1 0 5152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _396_
timestamp 1669390400
transform -1 0 19040 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _397_
timestamp 1669390400
transform -1 0 6384 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _398_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11760 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _399_
timestamp 1669390400
transform 1 0 12432 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _400_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6384 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _401_
timestamp 1669390400
transform 1 0 12432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _402_
timestamp 1669390400
transform 1 0 7952 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _403_
timestamp 1669390400
transform 1 0 8624 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _404_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 24976 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _405_
timestamp 1669390400
transform 1 0 14784 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _406_
timestamp 1669390400
transform 1 0 13552 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _407_
timestamp 1669390400
transform -1 0 14336 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _408_
timestamp 1669390400
transform -1 0 22960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _409_
timestamp 1669390400
transform -1 0 22960 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _410_
timestamp 1669390400
transform 1 0 18816 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _411_
timestamp 1669390400
transform -1 0 15232 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _412_
timestamp 1669390400
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _413_
timestamp 1669390400
transform 1 0 4480 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _414_
timestamp 1669390400
transform -1 0 25872 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _415_
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1669390400
transform -1 0 22848 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _417_
timestamp 1669390400
transform 1 0 5152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _418_
timestamp 1669390400
transform 1 0 9408 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _419_
timestamp 1669390400
transform 1 0 4480 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _420_
timestamp 1669390400
transform 1 0 3808 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _421_
timestamp 1669390400
transform -1 0 2352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _422_
timestamp 1669390400
transform 1 0 4144 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _423_
timestamp 1669390400
transform 1 0 1792 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _424_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 21056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _425_
timestamp 1669390400
transform -1 0 10080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _426_
timestamp 1669390400
transform -1 0 9184 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _427_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7840 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _428_
timestamp 1669390400
transform -1 0 2352 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _429_
timestamp 1669390400
transform 1 0 7504 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _430_
timestamp 1669390400
transform 1 0 9744 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _431_
timestamp 1669390400
transform -1 0 26880 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _432_
timestamp 1669390400
transform 1 0 18256 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _433_
timestamp 1669390400
transform 1 0 21504 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _434_
timestamp 1669390400
transform -1 0 18816 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _435_
timestamp 1669390400
transform -1 0 33040 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _436_
timestamp 1669390400
transform 1 0 14000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _437_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21728 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _438_
timestamp 1669390400
transform -1 0 30800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _439_
timestamp 1669390400
transform 1 0 25536 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _440_
timestamp 1669390400
transform 1 0 29456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _441_
timestamp 1669390400
transform -1 0 27664 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _442_
timestamp 1669390400
transform 1 0 24080 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _443_
timestamp 1669390400
transform 1 0 29456 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _444_
timestamp 1669390400
transform -1 0 28560 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _445_
timestamp 1669390400
transform 1 0 29456 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _446_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 28112 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _447_
timestamp 1669390400
transform -1 0 28000 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _448_
timestamp 1669390400
transform -1 0 30800 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _449_
timestamp 1669390400
transform -1 0 28784 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _450_
timestamp 1669390400
transform 1 0 29904 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _451_
timestamp 1669390400
transform -1 0 29008 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _452_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _453_
timestamp 1669390400
transform 1 0 8288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _454_
timestamp 1669390400
transform -1 0 33040 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _455_
timestamp 1669390400
transform 1 0 30912 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _456_
timestamp 1669390400
transform 1 0 30128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _457_
timestamp 1669390400
transform 1 0 33488 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _458_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 28112 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _459_
timestamp 1669390400
transform -1 0 30688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _460_
timestamp 1669390400
transform 1 0 31584 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _461_
timestamp 1669390400
transform 1 0 30800 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _462_
timestamp 1669390400
transform -1 0 31472 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _463_
timestamp 1669390400
transform 1 0 32368 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _464_
timestamp 1669390400
transform -1 0 34048 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _465_
timestamp 1669390400
transform -1 0 30464 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _466_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 32144 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _467_
timestamp 1669390400
transform -1 0 35840 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _468_
timestamp 1669390400
transform 1 0 33488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _469_
timestamp 1669390400
transform 1 0 32368 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _470_
timestamp 1669390400
transform 1 0 31808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _471_
timestamp 1669390400
transform -1 0 36400 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _472_
timestamp 1669390400
transform -1 0 31136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _473_
timestamp 1669390400
transform 1 0 36064 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _474_
timestamp 1669390400
transform -1 0 31136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _475_
timestamp 1669390400
transform 1 0 29008 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _476_
timestamp 1669390400
transform 1 0 32144 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _477_
timestamp 1669390400
transform -1 0 38864 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _478_
timestamp 1669390400
transform -1 0 38080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _479_
timestamp 1669390400
transform 1 0 31360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _480_
timestamp 1669390400
transform -1 0 36512 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _481_
timestamp 1669390400
transform 1 0 33488 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _482_
timestamp 1669390400
transform 1 0 34608 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _483_
timestamp 1669390400
transform -1 0 35616 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _484_
timestamp 1669390400
transform -1 0 36400 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _485_
timestamp 1669390400
transform -1 0 36512 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _486_
timestamp 1669390400
transform -1 0 39536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _487_
timestamp 1669390400
transform -1 0 37184 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _488_
timestamp 1669390400
transform -1 0 35616 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _489_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 39760 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _490_
timestamp 1669390400
transform 1 0 37520 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _491_
timestamp 1669390400
transform 1 0 37408 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _492_
timestamp 1669390400
transform -1 0 39424 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _493_
timestamp 1669390400
transform 1 0 37856 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _494_
timestamp 1669390400
transform -1 0 38304 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _495_
timestamp 1669390400
transform -1 0 39200 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _496_
timestamp 1669390400
transform -1 0 38864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _497_
timestamp 1669390400
transform -1 0 38304 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _498_
timestamp 1669390400
transform 1 0 8624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _499_
timestamp 1669390400
transform 1 0 6720 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _500_
timestamp 1669390400
transform 1 0 9632 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _501_
timestamp 1669390400
transform 1 0 9632 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _502_
timestamp 1669390400
transform 1 0 9632 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _503_
timestamp 1669390400
transform 1 0 6160 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _504_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7056 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _505_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6832 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _506_
timestamp 1669390400
transform 1 0 1792 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _507_
timestamp 1669390400
transform 1 0 2128 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _508_
timestamp 1669390400
transform 1 0 7840 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1669390400
transform -1 0 8736 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _510_
timestamp 1669390400
transform 1 0 7392 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _511_
timestamp 1669390400
transform 1 0 6048 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _512_
timestamp 1669390400
transform 1 0 2128 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _513_
timestamp 1669390400
transform -1 0 7728 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _514_
timestamp 1669390400
transform 1 0 6048 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _515_
timestamp 1669390400
transform 1 0 2352 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _516_
timestamp 1669390400
transform 1 0 2576 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _517_
timestamp 1669390400
transform 1 0 5040 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _518_
timestamp 1669390400
transform -1 0 8960 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _519_
timestamp 1669390400
transform -1 0 6832 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _520_
timestamp 1669390400
transform 1 0 3360 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _521_
timestamp 1669390400
transform -1 0 6720 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _522_
timestamp 1669390400
transform 1 0 6944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _523_
timestamp 1669390400
transform -1 0 6720 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _524_
timestamp 1669390400
transform 1 0 1680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _525_
timestamp 1669390400
transform 1 0 1680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _526_
timestamp 1669390400
transform 1 0 2576 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _527_
timestamp 1669390400
transform -1 0 8064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _528_
timestamp 1669390400
transform -1 0 8736 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _529_
timestamp 1669390400
transform 1 0 5040 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _530_
timestamp 1669390400
transform 1 0 5600 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _531_
timestamp 1669390400
transform 1 0 1792 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _532_
timestamp 1669390400
transform 1 0 3472 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _533_
timestamp 1669390400
transform 1 0 2576 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _534_
timestamp 1669390400
transform -1 0 3360 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _535_
timestamp 1669390400
transform 1 0 2352 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _536_
timestamp 1669390400
transform -1 0 4256 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _537_
timestamp 1669390400
transform 1 0 7056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _538_
timestamp 1669390400
transform 1 0 6608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _539_
timestamp 1669390400
transform 1 0 5600 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _540_
timestamp 1669390400
transform 1 0 3808 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _541_
timestamp 1669390400
transform -1 0 4144 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _542_
timestamp 1669390400
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _543_
timestamp 1669390400
transform 1 0 7056 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _544_
timestamp 1669390400
transform 1 0 2912 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _545_
timestamp 1669390400
transform 1 0 5264 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _546_
timestamp 1669390400
transform -1 0 6272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _547_
timestamp 1669390400
transform -1 0 6272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _548_
timestamp 1669390400
transform 1 0 8064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _549_
timestamp 1669390400
transform 1 0 7056 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _550_
timestamp 1669390400
transform 1 0 7840 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _551_
timestamp 1669390400
transform -1 0 9968 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _552_
timestamp 1669390400
transform 1 0 1680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _553_
timestamp 1669390400
transform 1 0 6832 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _554_
timestamp 1669390400
transform 1 0 4928 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _555_
timestamp 1669390400
transform -1 0 5600 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _556_
timestamp 1669390400
transform 1 0 3584 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _557_
timestamp 1669390400
transform 1 0 5600 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _558_
timestamp 1669390400
transform -1 0 7952 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _559_
timestamp 1669390400
transform 1 0 4144 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _560_
timestamp 1669390400
transform 1 0 6496 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _561_
timestamp 1669390400
transform 1 0 6944 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _562_
timestamp 1669390400
transform -1 0 10864 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _563_
timestamp 1669390400
transform -1 0 9184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _564_
timestamp 1669390400
transform 1 0 7952 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _565_
timestamp 1669390400
transform 1 0 4256 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _566_
timestamp 1669390400
transform 1 0 3360 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _567_
timestamp 1669390400
transform 1 0 6944 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _568_
timestamp 1669390400
transform 1 0 3360 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _569_
timestamp 1669390400
transform 1 0 4368 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _570_
timestamp 1669390400
transform 1 0 3696 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _571_
timestamp 1669390400
transform -1 0 6608 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _572_
timestamp 1669390400
transform 1 0 14448 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _573_
timestamp 1669390400
transform 1 0 15232 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _574_
timestamp 1669390400
transform 1 0 10080 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _575_
timestamp 1669390400
transform 1 0 9856 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _576_
timestamp 1669390400
transform 1 0 10976 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _577_
timestamp 1669390400
transform 1 0 13552 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _578_
timestamp 1669390400
transform -1 0 13776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _579_
timestamp 1669390400
transform 1 0 11760 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _580_
timestamp 1669390400
transform 1 0 12208 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _581_
timestamp 1669390400
transform 1 0 10192 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _582_
timestamp 1669390400
transform 1 0 9744 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _583_
timestamp 1669390400
transform 1 0 12544 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _584_
timestamp 1669390400
transform 1 0 10640 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _585_
timestamp 1669390400
transform 1 0 11424 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _586_
timestamp 1669390400
transform 1 0 14000 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _587_
timestamp 1669390400
transform 1 0 14560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _588_
timestamp 1669390400
transform 1 0 13440 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _589_
timestamp 1669390400
transform -1 0 14448 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _590_
timestamp 1669390400
transform 1 0 11200 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _591_
timestamp 1669390400
transform 1 0 13216 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _592_
timestamp 1669390400
transform 1 0 12544 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _593_
timestamp 1669390400
transform 1 0 14560 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _594_
timestamp 1669390400
transform -1 0 8400 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _595_
timestamp 1669390400
transform -1 0 8400 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _596_
timestamp 1669390400
transform 1 0 13104 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _597_
timestamp 1669390400
transform 1 0 14672 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _598_
timestamp 1669390400
transform 1 0 13888 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _599_
timestamp 1669390400
transform 1 0 14224 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _600_
timestamp 1669390400
transform -1 0 14784 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _601_
timestamp 1669390400
transform 1 0 12096 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _602_
timestamp 1669390400
transform 1 0 14560 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _603_
timestamp 1669390400
transform 1 0 12320 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _604_
timestamp 1669390400
transform -1 0 16016 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _605_
timestamp 1669390400
transform 1 0 15232 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _606_
timestamp 1669390400
transform -1 0 16352 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _607_
timestamp 1669390400
transform -1 0 16352 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _608_
timestamp 1669390400
transform -1 0 16240 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _609_
timestamp 1669390400
transform 1 0 13552 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _610_
timestamp 1669390400
transform 1 0 15792 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _611_
timestamp 1669390400
transform -1 0 16688 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _612_
timestamp 1669390400
transform 1 0 15680 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _613_
timestamp 1669390400
transform -1 0 18144 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _614_
timestamp 1669390400
transform 1 0 16576 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _615_
timestamp 1669390400
transform -1 0 16688 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _616_
timestamp 1669390400
transform 1 0 11088 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _617_
timestamp 1669390400
transform -1 0 11200 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _618_
timestamp 1669390400
transform 1 0 12544 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _619_
timestamp 1669390400
transform -1 0 16912 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _620_
timestamp 1669390400
transform 1 0 11536 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _621_
timestamp 1669390400
transform -1 0 16800 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _622_
timestamp 1669390400
transform -1 0 15904 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _623_
timestamp 1669390400
transform 1 0 16464 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _624_
timestamp 1669390400
transform 1 0 12096 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _625_
timestamp 1669390400
transform 1 0 17584 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _626_
timestamp 1669390400
transform 1 0 17584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1669390400
transform 1 0 4592 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _628_
timestamp 1669390400
transform 1 0 4592 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _629_
timestamp 1669390400
transform 1 0 15680 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _630_
timestamp 1669390400
transform 1 0 9632 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _631_
timestamp 1669390400
transform -1 0 18368 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _632_
timestamp 1669390400
transform -1 0 19488 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _633_
timestamp 1669390400
transform 1 0 16800 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _634_
timestamp 1669390400
transform 1 0 16688 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _635_
timestamp 1669390400
transform -1 0 17808 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _636_
timestamp 1669390400
transform 1 0 17808 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _637_
timestamp 1669390400
transform 1 0 15008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _638_
timestamp 1669390400
transform 1 0 18480 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1669390400
transform -1 0 25088 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _640_
timestamp 1669390400
transform 1 0 22960 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _641_
timestamp 1669390400
transform -1 0 22064 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _642_
timestamp 1669390400
transform 1 0 17584 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _643_
timestamp 1669390400
transform 1 0 19376 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _644_
timestamp 1669390400
transform 1 0 19264 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _645_
timestamp 1669390400
transform 1 0 20272 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _646_
timestamp 1669390400
transform 1 0 18592 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _647_
timestamp 1669390400
transform -1 0 21056 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _648_
timestamp 1669390400
transform 1 0 20160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _649_
timestamp 1669390400
transform -1 0 30464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _650_
timestamp 1669390400
transform 1 0 9072 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _651_
timestamp 1669390400
transform 1 0 10640 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _652_
timestamp 1669390400
transform -1 0 26880 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _653_
timestamp 1669390400
transform 1 0 21616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _654_
timestamp 1669390400
transform -1 0 21056 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _655_
timestamp 1669390400
transform 1 0 20272 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _656_
timestamp 1669390400
transform 1 0 18704 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1669390400
transform -1 0 24752 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _658_
timestamp 1669390400
transform 1 0 21728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _659_
timestamp 1669390400
transform -1 0 19600 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _660_
timestamp 1669390400
transform -1 0 18144 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _661_
timestamp 1669390400
transform 1 0 17584 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _662_
timestamp 1669390400
transform 1 0 16688 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _663_
timestamp 1669390400
transform -1 0 17584 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _664_
timestamp 1669390400
transform -1 0 18144 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _665_
timestamp 1669390400
transform 1 0 12544 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _666_
timestamp 1669390400
transform 1 0 18256 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _667_
timestamp 1669390400
transform 1 0 16576 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _668_
timestamp 1669390400
transform 1 0 17920 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1669390400
transform 1 0 17808 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _670_
timestamp 1669390400
transform 1 0 18592 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _671_
timestamp 1669390400
transform 1 0 19376 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _672_
timestamp 1669390400
transform 1 0 19600 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _673_
timestamp 1669390400
transform -1 0 19936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _674_
timestamp 1669390400
transform 1 0 18368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1669390400
transform 1 0 18368 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _676_
timestamp 1669390400
transform 1 0 18592 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _677_
timestamp 1669390400
transform -1 0 21952 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _678_
timestamp 1669390400
transform -1 0 22512 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1669390400
transform -1 0 20496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _680_
timestamp 1669390400
transform 1 0 19264 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _681_
timestamp 1669390400
transform -1 0 20720 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _682_
timestamp 1669390400
transform 1 0 20160 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _683_
timestamp 1669390400
transform -1 0 19712 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _684_
timestamp 1669390400
transform 1 0 20048 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _685_
timestamp 1669390400
transform 1 0 21504 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _686_
timestamp 1669390400
transform -1 0 23856 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _687_
timestamp 1669390400
transform -1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _688_
timestamp 1669390400
transform 1 0 19936 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _689_
timestamp 1669390400
transform 1 0 21392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _690_
timestamp 1669390400
transform -1 0 22400 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _691_
timestamp 1669390400
transform 1 0 24304 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _692_
timestamp 1669390400
transform -1 0 27664 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _693_
timestamp 1669390400
transform -1 0 26096 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _694_
timestamp 1669390400
transform -1 0 23968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _695_
timestamp 1669390400
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _696_
timestamp 1669390400
transform 1 0 24304 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _697_
timestamp 1669390400
transform 1 0 23184 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _698_
timestamp 1669390400
transform -1 0 24304 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _699_
timestamp 1669390400
transform 1 0 24192 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _700_
timestamp 1669390400
transform 1 0 25536 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1669390400
transform 1 0 27216 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _702_
timestamp 1669390400
transform -1 0 27104 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _703_
timestamp 1669390400
transform -1 0 28448 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _704_
timestamp 1669390400
transform 1 0 25984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _705_
timestamp 1669390400
transform -1 0 28896 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _706_
timestamp 1669390400
transform 1 0 26096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _707_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 23408 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1669390400
transform -1 0 22624 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _709_
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1669390400
transform 1 0 23744 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _711_
timestamp 1669390400
transform -1 0 28784 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _712_
timestamp 1669390400
transform 1 0 25872 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _713_
timestamp 1669390400
transform 1 0 28224 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1669390400
transform 1 0 29344 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _715_
timestamp 1669390400
transform 1 0 32368 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _716_
timestamp 1669390400
transform 1 0 31024 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _717_
timestamp 1669390400
transform 1 0 29792 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1669390400
transform 1 0 34496 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1669390400
transform 1 0 34496 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1669390400
transform 1 0 34608 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _721_
timestamp 1669390400
transform 1 0 33712 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _722_
timestamp 1669390400
transform 1 0 34496 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1669390400
transform -1 0 11536 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _724_
timestamp 1669390400
transform -1 0 6160 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _725_
timestamp 1669390400
transform 1 0 1680 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _726_
timestamp 1669390400
transform -1 0 4928 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _727_
timestamp 1669390400
transform -1 0 4928 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _728_
timestamp 1669390400
transform -1 0 4928 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _729_
timestamp 1669390400
transform -1 0 5040 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _730_
timestamp 1669390400
transform 1 0 7504 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _731_
timestamp 1669390400
transform -1 0 11872 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _732_
timestamp 1669390400
transform -1 0 12208 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _733_
timestamp 1669390400
transform -1 0 12768 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _734_
timestamp 1669390400
transform -1 0 15008 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _735_
timestamp 1669390400
transform 1 0 13776 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _736_
timestamp 1669390400
transform 1 0 16688 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _737_
timestamp 1669390400
transform 1 0 20608 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _738_
timestamp 1669390400
transform 1 0 21840 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _739_
timestamp 1669390400
transform 1 0 19376 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _740_
timestamp 1669390400
transform 1 0 22848 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _741_
timestamp 1669390400
transform 1 0 23184 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _742_
timestamp 1669390400
transform 1 0 26544 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _743_
timestamp 1669390400
transform 1 0 9744 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _744_
timestamp 1669390400
transform 1 0 10304 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18368 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform 1 0 22848 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform -1 0 28448 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input1 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16464 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 16464 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform -1 0 16912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform -1 0 19936 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 20832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform -1 0 23184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform 1 0 2576 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform 1 0 3360 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 5264 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 8064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform -1 0 9184 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform 1 0 7392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform 1 0 7280 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform 1 0 11984 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform 1 0 11200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform 1 0 1680 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38752 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 24416 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform -1 0 39536 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform -1 0 40320 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform -1 0 40320 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform 1 0 40544 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform -1 0 40320 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform -1 0 40320 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform -1 0 26768 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 26992 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform -1 0 28784 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform -1 0 31024 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 32480 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform 1 0 33040 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform 1 0 34832 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform -1 0 38528 0 1 3136
box -86 -86 1654 870
<< labels >>
flabel metal3 s 43200 21952 44000 22064 0 FreeSans 448 0 0 0 bs
port 0 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 clk
port 1 nsew signal input
flabel metal2 s 1120 0 1232 800 0 FreeSans 448 90 0 0 co[0]
port 2 nsew signal input
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 co[10]
port 3 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 co[11]
port 4 nsew signal input
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 co[12]
port 5 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 co[13]
port 6 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 co[14]
port 7 nsew signal input
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 co[15]
port 8 nsew signal input
flabel metal2 s 2464 0 2576 800 0 FreeSans 448 90 0 0 co[1]
port 9 nsew signal input
flabel metal2 s 3808 0 3920 800 0 FreeSans 448 90 0 0 co[2]
port 10 nsew signal input
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 co[3]
port 11 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 co[4]
port 12 nsew signal input
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 co[5]
port 13 nsew signal input
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 co[6]
port 14 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 co[7]
port 15 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 co[8]
port 16 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 co[9]
port 17 nsew signal input
flabel metal3 s 0 10976 800 11088 0 FreeSans 448 0 0 0 st
port 18 nsew signal input
flabel metal4 s 4448 3076 4768 40828 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 35168 3076 35488 40828 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 19808 3076 20128 40828 0 FreeSans 1280 90 0 0 vss
port 20 nsew ground bidirectional
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 x[0]
port 21 nsew signal tristate
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 x[10]
port 22 nsew signal tristate
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 x[11]
port 23 nsew signal tristate
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 x[12]
port 24 nsew signal tristate
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 x[13]
port 25 nsew signal tristate
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 x[14]
port 26 nsew signal tristate
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 x[15]
port 27 nsew signal tristate
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 x[1]
port 28 nsew signal tristate
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 x[2]
port 29 nsew signal tristate
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 x[3]
port 30 nsew signal tristate
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 x[4]
port 31 nsew signal tristate
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 x[5]
port 32 nsew signal tristate
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 x[6]
port 33 nsew signal tristate
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 x[7]
port 34 nsew signal tristate
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 x[8]
port 35 nsew signal tristate
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 x[9]
port 36 nsew signal tristate
rlabel metal1 21952 39984 21952 39984 0 vdd
rlabel metal1 21952 40768 21952 40768 0 vss
rlabel metal2 20328 5712 20328 5712 0 Datapath.i\[0\]
rlabel metal2 38808 10248 38808 10248 0 Datapath.i\[10\]
rlabel metal2 41944 6440 41944 6440 0 Datapath.i\[11\]
rlabel metal3 39984 5992 39984 5992 0 Datapath.i\[12\]
rlabel metal3 40264 7560 40264 7560 0 Datapath.i\[13\]
rlabel metal2 36792 11760 36792 11760 0 Datapath.i\[14\]
rlabel metal2 39032 9296 39032 9296 0 Datapath.i\[15\]
rlabel metal2 17640 4088 17640 4088 0 Datapath.i\[1\]
rlabel metal3 29736 15512 29736 15512 0 Datapath.i\[2\]
rlabel metal4 26824 12208 26824 12208 0 Datapath.i\[3\]
rlabel metal2 27776 15848 27776 15848 0 Datapath.i\[4\]
rlabel metal2 32256 15176 32256 15176 0 Datapath.i\[5\]
rlabel metal2 31696 11368 31696 11368 0 Datapath.i\[6\]
rlabel metal3 32144 10472 32144 10472 0 Datapath.i\[7\]
rlabel metal2 35448 9800 35448 9800 0 Datapath.i\[8\]
rlabel metal3 35224 8008 35224 8008 0 Datapath.i\[9\]
rlabel metal2 8456 5096 8456 5096 0 Datapath.k\[0\]
rlabel metal2 8568 21392 8568 21392 0 Datapath.k\[10\]
rlabel metal2 14896 17416 14896 17416 0 Datapath.k\[11\]
rlabel metal2 3192 22960 3192 22960 0 Datapath.k\[12\]
rlabel metal2 22568 19152 22568 19152 0 Datapath.k\[13\]
rlabel metal2 17640 22792 17640 22792 0 Datapath.k\[14\]
rlabel metal2 19656 18704 19656 18704 0 Datapath.k\[15\]
rlabel metal3 20888 17416 20888 17416 0 Datapath.k\[16\]
rlabel metal2 27160 15680 27160 15680 0 Datapath.k\[17\]
rlabel metal2 24528 12152 24528 12152 0 Datapath.k\[18\]
rlabel metal2 25816 11424 25816 11424 0 Datapath.k\[19\]
rlabel metal2 2408 16072 2408 16072 0 Datapath.k\[1\]
rlabel metal3 5096 9016 5096 9016 0 Datapath.k\[2\]
rlabel metal2 3080 22904 3080 22904 0 Datapath.k\[3\]
rlabel metal2 1904 8904 1904 8904 0 Datapath.k\[4\]
rlabel metal2 2688 20216 2688 20216 0 Datapath.k\[5\]
rlabel metal2 4760 20496 4760 20496 0 Datapath.k\[6\]
rlabel metal2 10024 15456 10024 15456 0 Datapath.k\[7\]
rlabel metal3 9128 19096 9128 19096 0 Datapath.k\[8\]
rlabel metal3 9352 15288 9352 15288 0 Datapath.k\[9\]
rlabel metal2 12656 9016 12656 9016 0 FSM.CS\[0\]
rlabel metal2 13384 4536 13384 4536 0 FSM.CS\[1\]
rlabel metal2 10696 7728 10696 7728 0 FSM.NS\[0\]
rlabel metal3 20720 22344 20720 22344 0 FSM.NS\[1\]
rlabel metal3 22120 5992 22120 5992 0 _000_
rlabel metal3 21952 4424 21952 4424 0 _001_
rlabel metal2 26488 4872 26488 4872 0 _002_
rlabel metal2 27832 5488 27832 5488 0 _003_
rlabel metal3 29064 8904 29064 8904 0 _004_
rlabel metal2 27384 10248 27384 10248 0 _005_
rlabel metal2 29176 8176 29176 8176 0 _006_
rlabel metal2 30240 9912 30240 9912 0 _007_
rlabel metal3 33544 9912 33544 9912 0 _008_
rlabel metal2 32032 6776 32032 6776 0 _009_
rlabel metal3 31192 5208 31192 5208 0 _010_
rlabel metal2 35392 4424 35392 4424 0 _011_
rlabel metal2 35392 5992 35392 5992 0 _012_
rlabel metal3 36624 7560 36624 7560 0 _013_
rlabel metal3 36120 11256 36120 11256 0 _014_
rlabel metal3 36512 9128 36512 9128 0 _015_
rlabel metal2 10584 5264 10584 5264 0 _016_
rlabel metal2 5880 3920 5880 3920 0 _017_
rlabel metal2 2632 5488 2632 5488 0 _018_
rlabel metal2 3920 7560 3920 7560 0 _019_
rlabel metal2 3976 9352 3976 9352 0 _020_
rlabel metal2 4312 11032 4312 11032 0 _021_
rlabel metal2 7336 13328 7336 13328 0 _022_
rlabel metal2 8456 15736 8456 15736 0 _023_
rlabel metal3 10584 13944 10584 13944 0 _024_
rlabel metal2 11704 17304 11704 17304 0 _025_
rlabel metal2 12544 11480 12544 11480 0 _026_
rlabel metal2 14056 10192 14056 10192 0 _027_
rlabel metal3 13720 4312 13720 4312 0 _028_
rlabel metal2 17640 6272 17640 6272 0 _029_
rlabel metal2 20552 7056 20552 7056 0 _030_
rlabel metal2 22008 8456 22008 8456 0 _031_
rlabel metal2 20272 12264 20272 12264 0 _032_
rlabel metal2 23800 14672 23800 14672 0 _033_
rlabel metal2 24136 10024 24136 10024 0 _034_
rlabel metal3 26376 12376 26376 12376 0 _035_
rlabel metal2 18536 17304 18536 17304 0 _036_
rlabel metal2 15736 19264 15736 19264 0 _037_
rlabel metal2 15736 6440 15736 6440 0 _038_
rlabel metal2 40880 6664 40880 6664 0 _039_
rlabel metal2 40936 3696 40936 3696 0 _040_
rlabel metal2 11032 5600 11032 5600 0 _041_
rlabel metal2 23968 15848 23968 15848 0 _042_
rlabel metal2 42168 9632 42168 9632 0 _043_
rlabel metal2 26208 15512 26208 15512 0 _044_
rlabel metal3 29680 15176 29680 15176 0 _045_
rlabel metal2 18312 20384 18312 20384 0 _046_
rlabel metal2 41608 9240 41608 9240 0 _047_
rlabel metal2 26824 6552 26824 6552 0 _048_
rlabel metal3 32928 4312 32928 4312 0 _049_
rlabel metal3 32480 8120 32480 8120 0 _050_
rlabel metal3 31472 8904 31472 8904 0 _051_
rlabel metal2 33992 11312 33992 11312 0 _052_
rlabel metal2 40320 8344 40320 8344 0 _053_
rlabel metal2 41832 4816 41832 4816 0 _054_
rlabel metal2 41944 4368 41944 4368 0 _055_
rlabel metal3 41216 7224 41216 7224 0 _056_
rlabel metal3 39872 8344 39872 8344 0 _057_
rlabel metal2 41608 6216 41608 6216 0 _058_
rlabel metal2 40096 5992 40096 5992 0 _059_
rlabel metal2 20888 17304 20888 17304 0 _060_
rlabel metal2 11816 21952 11816 21952 0 _061_
rlabel metal3 28952 15288 28952 15288 0 _062_
rlabel metal2 10080 23688 10080 23688 0 _063_
rlabel metal3 20608 15288 20608 15288 0 _064_
rlabel metal3 1904 18424 1904 18424 0 _065_
rlabel metal2 10472 7112 10472 7112 0 _066_
rlabel metal3 9072 2968 9072 2968 0 _067_
rlabel metal2 10248 3192 10248 3192 0 _068_
rlabel metal3 18200 21392 18200 21392 0 _069_
rlabel metal2 18088 4760 18088 4760 0 _070_
rlabel metal2 11928 5208 11928 5208 0 _071_
rlabel metal3 9520 4536 9520 4536 0 _072_
rlabel metal2 18984 20804 18984 20804 0 _073_
rlabel metal3 16464 2744 16464 2744 0 _074_
rlabel metal2 12712 17304 12712 17304 0 _075_
rlabel metal2 10360 17360 10360 17360 0 _076_
rlabel metal4 11704 13944 11704 13944 0 _077_
rlabel metal2 27664 15176 27664 15176 0 _078_
rlabel metal2 14728 18480 14728 18480 0 _079_
rlabel metal2 15400 17304 15400 17304 0 _080_
rlabel metal2 12600 14168 12600 14168 0 _081_
rlabel metal2 19152 12712 19152 12712 0 _082_
rlabel metal2 19040 12936 19040 12936 0 _083_
rlabel metal2 20608 15288 20608 15288 0 _084_
rlabel metal2 10248 9968 10248 9968 0 _085_
rlabel metal3 9240 17528 9240 17528 0 _086_
rlabel metal2 7784 11200 7784 11200 0 _087_
rlabel metal2 22568 12992 22568 12992 0 _088_
rlabel metal2 22680 17696 22680 17696 0 _089_
rlabel metal2 11424 22456 11424 22456 0 _090_
rlabel metal2 5432 9464 5432 9464 0 _091_
rlabel metal2 10136 9632 10136 9632 0 _092_
rlabel metal2 4760 16240 4760 16240 0 _093_
rlabel metal2 4088 19824 4088 19824 0 _094_
rlabel metal2 2968 21840 2968 21840 0 _095_
rlabel metal2 2296 19824 2296 19824 0 _096_
rlabel metal2 2408 21560 2408 21560 0 _097_
rlabel metal2 17976 18984 17976 18984 0 _098_
rlabel metal3 11424 19992 11424 19992 0 _099_
rlabel metal3 7448 24024 7448 24024 0 _100_
rlabel metal3 9520 7672 9520 7672 0 _101_
rlabel metal2 8904 22120 8904 22120 0 _102_
rlabel metal2 2744 22792 2744 22792 0 _103_
rlabel metal2 26712 11424 26712 11424 0 _104_
rlabel metal2 22344 8736 22344 8736 0 _105_
rlabel metal2 25816 16744 25816 16744 0 _106_
rlabel metal3 22792 17416 22792 17416 0 _107_
rlabel metal2 14392 5264 14392 5264 0 _108_
rlabel metal2 25704 6664 25704 6664 0 _109_
rlabel metal2 25816 9016 25816 9016 0 _110_
rlabel metal2 29792 12712 29792 12712 0 _111_
rlabel metal2 24808 5880 24808 5880 0 _112_
rlabel metal3 30632 15400 30632 15400 0 _113_
rlabel metal2 28056 9296 28056 9296 0 _114_
rlabel metal2 29960 7560 29960 7560 0 _115_
rlabel metal2 27720 8400 27720 8400 0 _116_
rlabel metal3 28840 5992 28840 5992 0 _117_
rlabel metal2 28672 9576 28672 9576 0 _118_
rlabel metal3 28000 9912 28000 9912 0 _119_
rlabel metal2 6496 11368 6496 11368 0 _120_
rlabel metal3 40600 9800 40600 9800 0 _121_
rlabel metal3 32088 8232 32088 8232 0 _122_
rlabel metal2 31192 8904 31192 8904 0 _123_
rlabel metal2 33656 8120 33656 8120 0 _124_
rlabel metal3 30632 13944 30632 13944 0 _125_
rlabel metal2 30408 8848 30408 8848 0 _126_
rlabel metal3 31248 11144 31248 11144 0 _127_
rlabel metal2 32648 11368 32648 11368 0 _128_
rlabel metal2 33544 10864 33544 10864 0 _129_
rlabel metal3 31696 9240 31696 9240 0 _130_
rlabel metal2 35560 7952 35560 7952 0 _131_
rlabel metal2 35560 9520 35560 9520 0 _132_
rlabel metal2 32592 7560 32592 7560 0 _133_
rlabel metal3 33880 5992 33880 5992 0 _134_
rlabel metal3 30128 5880 30128 5880 0 _135_
rlabel metal3 33768 12040 33768 12040 0 _136_
rlabel metal2 29288 6328 29288 6328 0 _137_
rlabel metal3 30744 5992 30744 5992 0 _138_
rlabel metal2 41944 9408 41944 9408 0 _139_
rlabel metal2 37912 5264 37912 5264 0 _140_
rlabel metal2 39704 10416 39704 10416 0 _141_
rlabel metal3 35056 5320 35056 5320 0 _142_
rlabel metal3 35224 6664 35224 6664 0 _143_
rlabel metal2 35000 7728 35000 7728 0 _144_
rlabel metal2 35672 6664 35672 6664 0 _145_
rlabel metal2 39368 8736 39368 8736 0 _146_
rlabel metal2 39200 9240 39200 9240 0 _147_
rlabel metal2 34888 6944 34888 6944 0 _148_
rlabel metal2 39256 11088 39256 11088 0 _149_
rlabel metal2 37800 7392 37800 7392 0 _150_
rlabel metal3 38192 11368 38192 11368 0 _151_
rlabel metal2 38248 10416 38248 10416 0 _152_
rlabel metal3 38192 9912 38192 9912 0 _153_
rlabel metal2 38136 9240 38136 9240 0 _154_
rlabel metal3 8120 7672 8120 7672 0 _155_
rlabel metal2 10248 5824 10248 5824 0 _156_
rlabel metal4 9912 20720 9912 20720 0 _157_
rlabel metal2 2968 13608 2968 13608 0 _158_
rlabel metal2 21896 18536 21896 18536 0 _159_
rlabel metal2 2744 5712 2744 5712 0 _160_
rlabel metal2 7896 24416 7896 24416 0 _161_
rlabel metal2 6048 24584 6048 24584 0 _162_
rlabel metal2 8288 17416 8288 17416 0 _163_
rlabel metal3 7448 11032 7448 11032 0 _164_
rlabel metal3 6664 17416 6664 17416 0 _165_
rlabel metal3 5040 3192 5040 3192 0 _166_
rlabel metal2 3304 24248 3304 24248 0 _167_
rlabel metal2 3192 21056 3192 21056 0 _168_
rlabel metal2 8344 8736 8344 8736 0 _169_
rlabel metal3 3220 15512 3220 15512 0 _170_
rlabel metal3 7280 11928 7280 11928 0 _171_
rlabel metal2 3976 8512 3976 8512 0 _172_
rlabel metal3 4872 8008 4872 8008 0 _173_
rlabel metal3 7000 9128 7000 9128 0 _174_
rlabel metal2 7224 9296 7224 9296 0 _175_
rlabel metal2 3192 19376 3192 19376 0 _176_
rlabel metal3 2464 8456 2464 8456 0 _177_
rlabel metal3 2464 9912 2464 9912 0 _178_
rlabel metal3 2968 17640 2968 17640 0 _179_
rlabel metal2 7336 10360 7336 10360 0 _180_
rlabel metal2 5208 10920 5208 10920 0 _181_
rlabel metal2 4088 10080 4088 10080 0 _182_
rlabel metal2 4200 9520 4200 9520 0 _183_
rlabel metal2 2520 12544 2520 12544 0 _184_
rlabel metal2 3024 17080 3024 17080 0 _185_
rlabel metal3 3024 12152 3024 12152 0 _186_
rlabel metal2 3864 12544 3864 12544 0 _187_
rlabel metal2 6160 21784 6160 21784 0 _188_
rlabel metal2 7448 11480 7448 11480 0 _189_
rlabel metal2 4424 10864 4424 10864 0 _190_
rlabel metal3 5320 10808 5320 10808 0 _191_
rlabel metal2 3752 12488 3752 12488 0 _192_
rlabel metal3 6048 10024 6048 10024 0 _193_
rlabel metal3 7728 13048 7728 13048 0 _194_
rlabel metal2 5096 15680 5096 15680 0 _195_
rlabel metal2 5768 13272 5768 13272 0 _196_
rlabel metal2 6048 13160 6048 13160 0 _197_
rlabel metal3 5992 12992 5992 12992 0 _198_
rlabel metal2 8456 12544 8456 12544 0 _199_
rlabel metal3 7448 15848 7448 15848 0 _200_
rlabel metal3 7784 12712 7784 12712 0 _201_
rlabel metal2 7560 12656 7560 12656 0 _202_
rlabel metal2 1960 12432 1960 12432 0 _203_
rlabel metal3 6440 15512 6440 15512 0 _204_
rlabel metal3 4424 16968 4424 16968 0 _205_
rlabel metal2 5992 16408 5992 16408 0 _206_
rlabel metal3 6944 16296 6944 16296 0 _207_
rlabel metal2 7560 16072 7560 16072 0 _208_
rlabel metal3 5600 15288 5600 15288 0 _209_
rlabel metal2 7168 15400 7168 15400 0 _210_
rlabel metal3 8064 15176 8064 15176 0 _211_
rlabel metal3 9072 15512 9072 15512 0 _212_
rlabel metal3 9520 16968 9520 16968 0 _213_
rlabel metal2 4872 16856 4872 16856 0 _214_
rlabel metal2 4536 12712 4536 12712 0 _215_
rlabel metal2 7448 14000 7448 14000 0 _216_
rlabel metal2 16184 15232 16184 15232 0 _217_
rlabel metal2 4648 12656 4648 12656 0 _218_
rlabel metal3 5040 15400 5040 15400 0 _219_
rlabel metal2 15176 16408 15176 16408 0 _220_
rlabel metal2 14952 15568 14952 15568 0 _221_
rlabel metal3 16464 15960 16464 15960 0 _222_
rlabel metal2 11256 16408 11256 16408 0 _223_
rlabel metal2 12712 15848 12712 15848 0 _224_
rlabel metal3 11704 15960 11704 15960 0 _225_
rlabel metal2 13944 17248 13944 17248 0 _226_
rlabel metal3 13160 15960 13160 15960 0 _227_
rlabel metal2 12264 15568 12264 15568 0 _228_
rlabel metal3 11424 15176 11424 15176 0 _229_
rlabel metal2 10472 12432 10472 12432 0 _230_
rlabel metal2 13832 16632 13832 16632 0 _231_
rlabel metal3 12152 15288 12152 15288 0 _232_
rlabel metal2 13384 16576 13384 16576 0 _233_
rlabel metal2 14616 16968 14616 16968 0 _234_
rlabel metal2 14840 16744 14840 16744 0 _235_
rlabel metal2 13720 16800 13720 16800 0 _236_
rlabel metal3 12712 16968 12712 16968 0 _237_
rlabel metal2 16408 15792 16408 15792 0 _238_
rlabel metal3 16632 15288 16632 15288 0 _239_
rlabel metal2 14168 14504 14168 14504 0 _240_
rlabel metal2 13384 13776 13384 13776 0 _241_
rlabel metal2 15568 18984 15568 18984 0 _242_
rlabel metal3 15680 14504 15680 14504 0 _243_
rlabel metal2 15400 13664 15400 13664 0 _244_
rlabel metal2 14392 14056 14392 14056 0 _245_
rlabel metal2 12712 12432 12712 12432 0 _246_
rlabel metal2 12936 9968 12936 9968 0 _247_
rlabel metal2 16184 18144 16184 18144 0 _248_
rlabel metal3 14336 13832 14336 13832 0 _249_
rlabel metal2 15512 12208 15512 12208 0 _250_
rlabel metal2 15736 11032 15736 11032 0 _251_
rlabel metal2 15960 12152 15960 12152 0 _252_
rlabel metal2 15624 10584 15624 10584 0 _253_
rlabel metal2 15288 7280 15288 7280 0 _254_
rlabel metal2 16520 15736 16520 15736 0 _255_
rlabel metal2 16296 15568 16296 15568 0 _256_
rlabel metal3 16856 11368 16856 11368 0 _257_
rlabel metal2 17640 15204 17640 15204 0 _258_
rlabel metal3 17080 11144 17080 11144 0 _259_
rlabel metal2 16856 17808 16856 17808 0 _260_
rlabel metal2 16296 9800 16296 9800 0 _261_
rlabel metal3 16912 18984 16912 18984 0 _262_
rlabel metal2 15848 19376 15848 19376 0 _263_
rlabel metal2 15736 9240 15736 9240 0 _264_
rlabel metal2 16072 17192 16072 17192 0 _265_
rlabel metal3 16072 9016 16072 9016 0 _266_
rlabel metal2 15400 8288 15400 8288 0 _267_
rlabel metal3 14896 6440 14896 6440 0 _268_
rlabel metal2 18032 16632 18032 16632 0 _269_
rlabel metal3 17304 9240 17304 9240 0 _270_
rlabel metal3 2240 23576 2240 23576 0 _271_
rlabel metal2 16968 18928 16968 18928 0 _272_
rlabel metal3 17080 7672 17080 7672 0 _273_
rlabel metal3 17976 20496 17976 20496 0 _274_
rlabel metal2 17416 7840 17416 7840 0 _275_
rlabel metal2 17640 8064 17640 8064 0 _276_
rlabel metal2 17192 10584 17192 10584 0 _277_
rlabel metal3 20216 11144 20216 11144 0 _278_
rlabel metal3 15512 10920 15512 10920 0 _279_
rlabel metal2 19656 10976 19656 10976 0 _280_
rlabel metal2 19656 9800 19656 9800 0 _281_
rlabel metal2 24528 11368 24528 11368 0 _282_
rlabel metal3 20160 9240 20160 9240 0 _283_
rlabel metal3 20496 11368 20496 11368 0 _284_
rlabel metal3 18704 9688 18704 9688 0 _285_
rlabel metal2 20440 9464 20440 9464 0 _286_
rlabel metal2 20272 8232 20272 8232 0 _287_
rlabel metal2 20440 7504 20440 7504 0 _288_
rlabel metal2 20216 7000 20216 7000 0 _289_
rlabel metal3 21280 9576 21280 9576 0 _290_
rlabel metal2 25648 5880 25648 5880 0 _291_
rlabel metal2 10808 9240 10808 9240 0 _292_
rlabel metal2 19208 16912 19208 16912 0 _293_
rlabel metal2 22456 9072 22456 9072 0 _294_
rlabel metal2 21896 9968 21896 9968 0 _295_
rlabel metal2 20776 10024 20776 10024 0 _296_
rlabel metal2 22232 8344 22232 8344 0 _297_
rlabel metal2 19880 8064 19880 8064 0 _298_
rlabel metal3 23464 7672 23464 7672 0 _299_
rlabel metal2 18648 9856 18648 9856 0 _300_
rlabel metal2 17696 10808 17696 10808 0 _301_
rlabel metal2 17864 13496 17864 13496 0 _302_
rlabel metal2 17416 15344 17416 15344 0 _303_
rlabel metal3 18760 15344 18760 15344 0 _304_
rlabel metal2 17640 12600 17640 12600 0 _305_
rlabel metal2 18872 9688 18872 9688 0 _306_
rlabel metal2 18536 10024 18536 10024 0 _307_
rlabel metal2 18088 14280 18088 14280 0 _308_
rlabel metal2 19600 17080 19600 17080 0 _309_
rlabel metal3 18872 13496 18872 13496 0 _310_
rlabel metal3 19264 15960 19264 15960 0 _311_
rlabel metal2 19768 15456 19768 15456 0 _312_
rlabel metal2 21336 15680 21336 15680 0 _313_
rlabel metal2 19208 15232 19208 15232 0 _314_
rlabel metal3 19208 15848 19208 15848 0 _315_
rlabel metal3 18984 15512 18984 15512 0 _316_
rlabel metal2 21448 16520 21448 16520 0 _317_
rlabel metal3 20664 12936 20664 12936 0 _318_
rlabel metal2 21896 11648 21896 11648 0 _319_
rlabel metal2 20776 15680 20776 15680 0 _320_
rlabel metal2 20216 14504 20216 14504 0 _321_
rlabel metal3 21504 15512 21504 15512 0 _322_
rlabel metal3 19824 14728 19824 14728 0 _323_
rlabel metal2 21560 16352 21560 16352 0 _324_
rlabel metal3 22512 15400 22512 15400 0 _325_
rlabel metal2 23352 12096 23352 12096 0 _326_
rlabel metal3 21448 14280 21448 14280 0 _327_
rlabel metal2 21672 14224 21672 14224 0 _328_
rlabel metal2 23352 13888 23352 13888 0 _329_
rlabel metal3 25424 12376 25424 12376 0 _330_
rlabel metal2 25984 13720 25984 13720 0 _331_
rlabel metal2 25536 12376 25536 12376 0 _332_
rlabel metal2 23576 13776 23576 13776 0 _333_
rlabel metal2 23800 12936 23800 12936 0 _334_
rlabel metal3 23968 13496 23968 13496 0 _335_
rlabel metal2 24584 10864 24584 10864 0 _336_
rlabel metal2 24248 10808 24248 10808 0 _337_
rlabel metal2 27384 12096 27384 12096 0 _338_
rlabel metal2 26712 13608 26712 13608 0 _339_
rlabel metal2 26376 14112 26376 14112 0 _340_
rlabel metal2 27944 13328 27944 13328 0 _341_
rlabel metal2 26264 13272 26264 13272 0 _342_
rlabel metal2 28392 11704 28392 11704 0 _343_
rlabel metal2 40040 22120 40040 22120 0 bs
rlabel metal3 854 32984 854 32984 0 clk
rlabel metal2 17640 19152 17640 19152 0 clknet_0_clk
rlabel metal3 20328 22120 20328 22120 0 clknet_2_0__leaf_clk
rlabel metal2 5656 21168 5656 21168 0 clknet_2_1__leaf_clk
rlabel metal2 29512 16464 29512 16464 0 clknet_2_2__leaf_clk
rlabel metal2 23520 9800 23520 9800 0 clknet_2_3__leaf_clk
rlabel metal2 1176 1638 1176 1638 0 co[0]
rlabel metal3 15680 21896 15680 21896 0 co[10]
rlabel metal2 42392 4760 42392 4760 0 co[11]
rlabel metal2 17304 1806 17304 1806 0 co[12]
rlabel metal2 19096 728 19096 728 0 co[13]
rlabel metal2 19992 1862 19992 1862 0 co[14]
rlabel metal3 22960 3416 22960 3416 0 co[15]
rlabel metal2 2744 2968 2744 2968 0 co[1]
rlabel metal3 23296 2632 23296 2632 0 co[2]
rlabel metal2 1288 14168 1288 14168 0 co[3]
rlabel metal2 1624 14336 1624 14336 0 co[4]
rlabel metal2 8904 6104 8904 6104 0 co[5]
rlabel metal3 5712 20328 5712 20328 0 co[6]
rlabel metal2 10584 2030 10584 2030 0 co[7]
rlabel metal3 12880 23576 12880 23576 0 co[8]
rlabel metal3 18592 21448 18592 21448 0 co[9]
rlabel metal3 11536 24024 11536 24024 0 net1
rlabel metal3 6384 7336 6384 7336 0 net10
rlabel metal2 6216 7504 6216 7504 0 net11
rlabel metal2 6776 21280 6776 21280 0 net12
rlabel metal2 1848 22512 1848 22512 0 net13
rlabel metal3 10472 3752 10472 3752 0 net14
rlabel metal3 17388 20664 17388 20664 0 net15
rlabel metal2 14056 4872 14056 4872 0 net16
rlabel metal2 3416 10976 3416 10976 0 net17
rlabel metal3 39984 8232 39984 8232 0 net18
rlabel metal2 23968 3752 23968 3752 0 net19
rlabel metal2 14784 5768 14784 5768 0 net2
rlabel metal2 39368 4368 39368 4368 0 net20
rlabel metal3 40880 3528 40880 3528 0 net21
rlabel metal2 39928 5376 39928 5376 0 net22
rlabel metal3 40096 5096 40096 5096 0 net23
rlabel metal2 41720 6384 41720 6384 0 net24
rlabel metal2 40264 6776 40264 6776 0 net25
rlabel metal2 27608 16968 27608 16968 0 net26
rlabel metal2 26936 16296 26936 16296 0 net27
rlabel metal2 28504 4816 28504 4816 0 net28
rlabel metal2 29512 6328 29512 6328 0 net29
rlabel metal2 16072 5880 16072 5880 0 net3
rlabel metal2 30856 4368 30856 4368 0 net30
rlabel metal2 32312 4704 32312 4704 0 net31
rlabel metal2 33152 3528 33152 3528 0 net32
rlabel metal2 35000 3808 35000 3808 0 net33
rlabel metal2 38360 3808 38360 3808 0 net34
rlabel metal3 16016 3640 16016 3640 0 net4
rlabel metal2 18536 6160 18536 6160 0 net5
rlabel metal2 18704 4312 18704 4312 0 net6
rlabel metal2 18760 4032 18760 4032 0 net7
rlabel via1 5768 19432 5768 19432 0 net8
rlabel metal2 5768 5880 5768 5880 0 net9
rlabel metal3 1302 11032 1302 11032 0 st
rlabel metal2 22680 2058 22680 2058 0 x[0]
rlabel metal3 37184 4200 37184 4200 0 x[10]
rlabel metal2 37464 2086 37464 2086 0 x[11]
rlabel metal2 38808 2870 38808 2870 0 x[12]
rlabel metal2 40152 1638 40152 1638 0 x[13]
rlabel metal2 41496 2198 41496 2198 0 x[14]
rlabel metal2 42840 2310 42840 2310 0 x[15]
rlabel metal3 24752 3416 24752 3416 0 x[1]
rlabel metal2 25368 2198 25368 2198 0 x[2]
rlabel metal2 26712 2870 26712 2870 0 x[3]
rlabel metal3 29008 3640 29008 3640 0 x[4]
rlabel metal2 29400 854 29400 854 0 x[5]
rlabel metal2 30744 2058 30744 2058 0 x[6]
rlabel metal2 32088 1246 32088 1246 0 x[7]
rlabel metal3 34552 3528 34552 3528 0 x[8]
rlabel metal3 36008 3416 36008 3416 0 x[9]
<< properties >>
string FIXED_BBOX 0 0 44000 44000
<< end >>
