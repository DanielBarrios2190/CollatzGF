// This is the unpowered netlist.
module collatz (bs,
    clk,
    st,
    co,
    x);
 output bs;
 input clk;
 input st;
 input [15:0] co;
 output [15:0] x;

 wire \Datapath.i[0] ;
 wire \Datapath.i[10] ;
 wire \Datapath.i[11] ;
 wire \Datapath.i[12] ;
 wire \Datapath.i[13] ;
 wire \Datapath.i[14] ;
 wire \Datapath.i[15] ;
 wire \Datapath.i[1] ;
 wire \Datapath.i[2] ;
 wire \Datapath.i[3] ;
 wire \Datapath.i[4] ;
 wire \Datapath.i[5] ;
 wire \Datapath.i[6] ;
 wire \Datapath.i[7] ;
 wire \Datapath.i[8] ;
 wire \Datapath.i[9] ;
 wire \Datapath.k[0] ;
 wire \Datapath.k[10] ;
 wire \Datapath.k[11] ;
 wire \Datapath.k[12] ;
 wire \Datapath.k[13] ;
 wire \Datapath.k[14] ;
 wire \Datapath.k[15] ;
 wire \Datapath.k[16] ;
 wire \Datapath.k[17] ;
 wire \Datapath.k[18] ;
 wire \Datapath.k[19] ;
 wire \Datapath.k[1] ;
 wire \Datapath.k[2] ;
 wire \Datapath.k[3] ;
 wire \Datapath.k[4] ;
 wire \Datapath.k[5] ;
 wire \Datapath.k[6] ;
 wire \Datapath.k[7] ;
 wire \Datapath.k[8] ;
 wire \Datapath.k[9] ;
 wire \FSM.CS[0] ;
 wire \FSM.CS[1] ;
 wire \FSM.NS[0] ;
 wire \FSM.NS[1] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__buf_4 _246_ (.I(\FSM.CS[0] ),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _247_ (.A1(_036_),
    .A2(\FSM.CS[1] ),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _248_ (.I(_037_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _249_ (.A1(\Datapath.i[0] ),
    .A2(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _250_ (.I(_038_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _251_ (.I(_037_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _252_ (.A1(\Datapath.i[1] ),
    .A2(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _253_ (.I(_040_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _254_ (.A1(\Datapath.i[2] ),
    .A2(_039_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _255_ (.I(_041_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _256_ (.A1(\Datapath.i[3] ),
    .A2(_039_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _257_ (.I(_042_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _258_ (.A1(\Datapath.i[4] ),
    .A2(_039_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _259_ (.I(_043_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _260_ (.A1(\Datapath.i[5] ),
    .A2(_039_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(_044_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _262_ (.A1(\Datapath.i[6] ),
    .A2(_039_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(_045_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _264_ (.A1(\Datapath.i[7] ),
    .A2(_039_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _265_ (.I(_046_),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _266_ (.A1(\Datapath.i[8] ),
    .A2(_039_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(_047_),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _268_ (.A1(\Datapath.i[9] ),
    .A2(_039_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(_048_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _270_ (.A1(\Datapath.i[10] ),
    .A2(_039_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _271_ (.I(_049_),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _272_ (.A1(\Datapath.i[11] ),
    .A2(_039_),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _273_ (.I(_050_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _274_ (.A1(\Datapath.i[12] ),
    .A2(_039_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _275_ (.I(_051_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _276_ (.A1(\Datapath.i[13] ),
    .A2(_039_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _277_ (.I(_052_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _278_ (.A1(\Datapath.i[14] ),
    .A2(_039_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _279_ (.I(_053_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _280_ (.A1(\Datapath.i[15] ),
    .A2(_037_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _281_ (.I(_054_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _282_ (.I(\FSM.CS[1] ),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _283_ (.A1(_036_),
    .A2(\Datapath.k[1] ),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _284_ (.A1(_055_),
    .A2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _285_ (.I(_036_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _286_ (.I(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _287_ (.A1(_058_),
    .A2(\FSM.CS[1] ),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _288_ (.I(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _289_ (.I(net1),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _290_ (.A1(_059_),
    .A2(net17),
    .B1(_061_),
    .B2(_062_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _291_ (.A1(_057_),
    .A2(_063_),
    .ZN(\FSM.NS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _292_ (.A1(net11),
    .A2(net12),
    .A3(net13),
    .A4(net14),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _293_ (.A1(_062_),
    .A2(net8),
    .A3(net9),
    .A4(net10),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _294_ (.A1(net15),
    .A2(net16),
    .A3(net2),
    .A4(net3),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _295_ (.A1(net4),
    .A2(net5),
    .A3(net6),
    .A4(net7),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _296_ (.A1(_064_),
    .A2(_065_),
    .A3(_066_),
    .A4(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _297_ (.A1(\Datapath.k[17] ),
    .A2(\Datapath.k[16] ),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _298_ (.I(\Datapath.k[9] ),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _299_ (.A1(\Datapath.k[13] ),
    .A2(\Datapath.k[12] ),
    .A3(_070_),
    .A4(\Datapath.k[8] ),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _300_ (.A1(\Datapath.k[3] ),
    .A2(\Datapath.k[2] ),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _301_ (.I(\Datapath.k[4] ),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _302_ (.A1(\Datapath.k[11] ),
    .A2(\Datapath.k[10] ),
    .A3(\Datapath.k[5] ),
    .A4(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _303_ (.A1(\Datapath.k[7] ),
    .A2(\Datapath.k[6] ),
    .A3(_072_),
    .A4(_074_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _304_ (.A1(\Datapath.k[19] ),
    .A2(\Datapath.k[18] ),
    .A3(\Datapath.k[15] ),
    .A4(\Datapath.k[14] ),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _305_ (.A1(\Datapath.k[0] ),
    .A2(_056_),
    .A3(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _306_ (.A1(_069_),
    .A2(_071_),
    .A3(_075_),
    .A4(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _307_ (.A1(_061_),
    .A2(_068_),
    .B1(_078_),
    .B2(_055_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _308_ (.I(_079_),
    .ZN(\FSM.NS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _309_ (.I(\FSM.CS[1] ),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _310_ (.A1(\Datapath.i[0] ),
    .A2(_080_),
    .B(_038_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _311_ (.A1(\Datapath.i[1] ),
    .A2(\Datapath.i[0] ),
    .A3(_055_),
    .Z(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _312_ (.A1(_036_),
    .A2(_080_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _313_ (.A1(\Datapath.i[0] ),
    .A2(_055_),
    .B1(_082_),
    .B2(\Datapath.i[1] ),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _314_ (.A1(_081_),
    .A2(_083_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _315_ (.A1(\Datapath.i[2] ),
    .A2(_081_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _316_ (.A1(\Datapath.i[2] ),
    .A2(\Datapath.i[1] ),
    .A3(\Datapath.i[0] ),
    .A4(\FSM.CS[1] ),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _317_ (.A1(_061_),
    .A2(_084_),
    .A3(_085_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _318_ (.A1(\Datapath.i[3] ),
    .A2(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _319_ (.A1(\Datapath.i[3] ),
    .A2(_085_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _320_ (.A1(_061_),
    .A2(_086_),
    .A3(_087_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _321_ (.A1(\Datapath.i[4] ),
    .A2(_087_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _322_ (.A1(\Datapath.i[4] ),
    .A2(_087_),
    .B(_082_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _323_ (.A1(_088_),
    .A2(_089_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _324_ (.A1(\Datapath.i[5] ),
    .A2(_088_),
    .B(_060_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _325_ (.A1(\Datapath.i[5] ),
    .A2(_088_),
    .B(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _326_ (.I(_091_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _327_ (.A1(\Datapath.i[5] ),
    .A2(_088_),
    .B(\Datapath.i[6] ),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _328_ (.A1(\Datapath.i[6] ),
    .A2(\Datapath.i[5] ),
    .A3(\Datapath.i[4] ),
    .A4(_087_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _329_ (.A1(_061_),
    .A2(_092_),
    .A3(_093_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _330_ (.A1(\Datapath.i[7] ),
    .A2(_093_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _331_ (.A1(\Datapath.i[7] ),
    .A2(_093_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _332_ (.A1(_061_),
    .A2(_094_),
    .A3(_095_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _333_ (.A1(\Datapath.i[8] ),
    .A2(\Datapath.i[7] ),
    .A3(_093_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _334_ (.A1(\Datapath.i[8] ),
    .A2(_095_),
    .B(_082_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _335_ (.A1(_096_),
    .A2(_097_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _336_ (.A1(\Datapath.i[9] ),
    .A2(_096_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _337_ (.A1(\Datapath.i[9] ),
    .A2(_096_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _338_ (.A1(_061_),
    .A2(_098_),
    .A3(_099_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _339_ (.A1(\Datapath.i[10] ),
    .A2(_099_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _340_ (.A1(\Datapath.i[10] ),
    .A2(_099_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _341_ (.A1(_061_),
    .A2(_100_),
    .A3(_101_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _342_ (.A1(\Datapath.i[11] ),
    .A2(_101_),
    .B(_060_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _343_ (.A1(\Datapath.i[11] ),
    .A2(_101_),
    .B(_102_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _344_ (.I(_103_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _345_ (.A1(\Datapath.i[11] ),
    .A2(_101_),
    .B(\Datapath.i[12] ),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _346_ (.A1(\Datapath.i[12] ),
    .A2(\Datapath.i[11] ),
    .A3(_101_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _347_ (.A1(_061_),
    .A2(_104_),
    .A3(_105_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _348_ (.A1(\Datapath.i[13] ),
    .A2(_105_),
    .B(_060_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _349_ (.A1(\Datapath.i[13] ),
    .A2(_105_),
    .B(_106_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _350_ (.I(_107_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _351_ (.A1(\Datapath.i[13] ),
    .A2(_105_),
    .B(\Datapath.i[14] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _352_ (.A1(\Datapath.i[14] ),
    .A2(\Datapath.i[13] ),
    .A3(_105_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _353_ (.A1(_061_),
    .A2(_108_),
    .A3(_109_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _354_ (.A1(\Datapath.i[15] ),
    .A2(_109_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _355_ (.A1(_082_),
    .A2(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _356_ (.I(_111_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _357_ (.A1(_036_),
    .A2(\Datapath.k[0] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _358_ (.A1(_057_),
    .A2(_112_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _359_ (.A1(_062_),
    .A2(_061_),
    .B1(_112_),
    .B2(_080_),
    .C(_113_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _360_ (.I(\Datapath.k[2] ),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _361_ (.A1(_036_),
    .A2(_055_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _362_ (.A1(_059_),
    .A2(\Datapath.k[1] ),
    .B1(net8),
    .B2(_061_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _363_ (.A1(_114_),
    .A2(_115_),
    .B(_116_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _364_ (.A1(\Datapath.k[2] ),
    .A2(\Datapath.k[1] ),
    .A3(\Datapath.k[0] ),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _365_ (.A1(_036_),
    .A2(_117_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _366_ (.A1(_055_),
    .A2(net9),
    .B1(_115_),
    .B2(\Datapath.k[3] ),
    .C(net18),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _367_ (.A1(_114_),
    .A2(net18),
    .B1(_118_),
    .B2(_119_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _368_ (.A1(\Datapath.k[3] ),
    .A2(net18),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _369_ (.I(\Datapath.k[0] ),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _370_ (.A1(\Datapath.k[2] ),
    .A2(\Datapath.k[1] ),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _371_ (.A1(\Datapath.k[2] ),
    .A2(\Datapath.k[1] ),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _372_ (.A1(_121_),
    .A2(_122_),
    .B(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _373_ (.A1(\Datapath.k[3] ),
    .A2(\Datapath.k[2] ),
    .A3(_124_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _374_ (.I0(_073_),
    .I1(_125_),
    .S(_059_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _375_ (.A1(_080_),
    .A2(net10),
    .B1(_082_),
    .B2(_126_),
    .C(_037_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _376_ (.A1(_120_),
    .A2(_127_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _377_ (.A1(_059_),
    .A2(_055_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _378_ (.A1(_073_),
    .A2(\Datapath.k[3] ),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _379_ (.A1(\Datapath.k[3] ),
    .A2(\Datapath.k[2] ),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _380_ (.A1(_121_),
    .A2(_122_),
    .B(_130_),
    .C(_123_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _381_ (.A1(_072_),
    .A2(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _382_ (.A1(_129_),
    .A2(_132_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _383_ (.A1(_128_),
    .A2(_133_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _384_ (.A1(_073_),
    .A2(net18),
    .B1(_082_),
    .B2(net11),
    .C1(_115_),
    .C2(\Datapath.k[5] ),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _385_ (.A1(_134_),
    .A2(_135_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _386_ (.A1(\Datapath.k[5] ),
    .A2(_073_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _387_ (.A1(_129_),
    .A2(_132_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _388_ (.A1(_073_),
    .A2(\Datapath.k[3] ),
    .B(_137_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _389_ (.A1(_136_),
    .A2(_138_),
    .Z(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _390_ (.A1(_036_),
    .A2(_139_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _391_ (.A1(_059_),
    .A2(\Datapath.k[6] ),
    .B(_055_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _392_ (.A1(\Datapath.k[5] ),
    .A2(_037_),
    .B1(_061_),
    .B2(net12),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _393_ (.A1(_140_),
    .A2(_141_),
    .B(_142_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _394_ (.A1(\Datapath.k[6] ),
    .A2(\Datapath.k[5] ),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _395_ (.A1(_073_),
    .A2(\Datapath.k[3] ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _396_ (.A1(\Datapath.k[5] ),
    .A2(_073_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _397_ (.A1(_144_),
    .A2(_145_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _398_ (.A1(\Datapath.k[5] ),
    .A2(_073_),
    .B1(_137_),
    .B2(_146_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _399_ (.A1(_143_),
    .A2(_147_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _400_ (.A1(_036_),
    .A2(_148_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _401_ (.A1(_055_),
    .A2(net13),
    .B1(_115_),
    .B2(\Datapath.k[7] ),
    .C(net18),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _402_ (.A1(\Datapath.k[6] ),
    .A2(_037_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _403_ (.A1(_149_),
    .A2(_150_),
    .B(_151_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _404_ (.A1(\Datapath.k[7] ),
    .A2(\Datapath.k[6] ),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _405_ (.A1(\Datapath.k[6] ),
    .A2(\Datapath.k[5] ),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _406_ (.A1(_143_),
    .A2(_147_),
    .B(_153_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _407_ (.A1(_152_),
    .A2(_154_),
    .B(_059_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _408_ (.A1(_152_),
    .A2(_154_),
    .B(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _409_ (.A1(_059_),
    .A2(\Datapath.k[8] ),
    .B(_055_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _410_ (.A1(\Datapath.k[7] ),
    .A2(_037_),
    .B1(_060_),
    .B2(net14),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _411_ (.A1(_156_),
    .A2(_157_),
    .B(_158_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _412_ (.A1(_036_),
    .A2(_080_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _413_ (.A1(_129_),
    .A2(_136_),
    .A3(_143_),
    .A4(_152_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _414_ (.A1(_072_),
    .A2(_131_),
    .A3(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _415_ (.A1(_144_),
    .A2(_145_),
    .B(_143_),
    .C(_152_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _416_ (.A1(\Datapath.k[7] ),
    .A2(\Datapath.k[6] ),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _417_ (.A1(_153_),
    .A2(_163_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _418_ (.A1(_161_),
    .A2(_162_),
    .A3(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _419_ (.A1(\Datapath.k[8] ),
    .A2(\Datapath.k[7] ),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _420_ (.A1(_165_),
    .A2(_166_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _421_ (.A1(\Datapath.k[8] ),
    .A2(net18),
    .B1(_082_),
    .B2(net15),
    .C1(_115_),
    .C2(_070_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _422_ (.A1(_159_),
    .A2(_167_),
    .B(_168_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _423_ (.A1(_059_),
    .A2(\Datapath.k[10] ),
    .B(_055_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _424_ (.A1(_070_),
    .A2(\Datapath.k[8] ),
    .Z(_170_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _425_ (.I(_166_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _426_ (.A1(\Datapath.k[8] ),
    .A2(\Datapath.k[7] ),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _427_ (.A1(_165_),
    .A2(_171_),
    .B(_172_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _428_ (.A1(_170_),
    .A2(_173_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _429_ (.A1(_036_),
    .A2(_174_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _430_ (.A1(_070_),
    .A2(_037_),
    .B1(_060_),
    .B2(net16),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _431_ (.A1(_169_),
    .A2(_175_),
    .B(_176_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _432_ (.A1(\Datapath.k[10] ),
    .A2(_070_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _433_ (.A1(_165_),
    .A2(_171_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _434_ (.A1(_070_),
    .A2(\Datapath.k[8] ),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _435_ (.A1(_172_),
    .A2(_179_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _436_ (.A1(_070_),
    .A2(\Datapath.k[8] ),
    .B1(_178_),
    .B2(_180_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _437_ (.A1(_177_),
    .A2(_181_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _438_ (.I0(\Datapath.k[11] ),
    .I1(net2),
    .I2(_182_),
    .I3(\Datapath.k[10] ),
    .S0(_080_),
    .S1(_059_),
    .Z(_183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _439_ (.I(_183_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _440_ (.A1(\Datapath.k[11] ),
    .A2(\Datapath.k[10] ),
    .Z(_184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _441_ (.A1(\Datapath.k[10] ),
    .A2(_070_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _442_ (.A1(\Datapath.k[10] ),
    .A2(_070_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _443_ (.A1(_185_),
    .A2(_181_),
    .B(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _444_ (.A1(_184_),
    .A2(_187_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _445_ (.A1(_036_),
    .A2(_188_),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _446_ (.A1(_059_),
    .A2(\Datapath.k[12] ),
    .B(_055_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _447_ (.A1(\Datapath.k[11] ),
    .A2(_037_),
    .B1(_060_),
    .B2(net3),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _448_ (.A1(_189_),
    .A2(_190_),
    .B(_191_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _449_ (.A1(_166_),
    .A2(_170_),
    .A3(_177_),
    .A4(_184_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _450_ (.A1(_161_),
    .A2(_162_),
    .A3(_164_),
    .B(_192_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _451_ (.A1(\Datapath.k[11] ),
    .A2(\Datapath.k[10] ),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _452_ (.A1(_177_),
    .A2(_180_),
    .A3(_184_),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _453_ (.A1(_186_),
    .A2(_194_),
    .A3(_195_),
    .Z(_196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _454_ (.A1(_193_),
    .A2(_196_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _455_ (.A1(\Datapath.k[12] ),
    .A2(\Datapath.k[11] ),
    .Z(_198_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _456_ (.A1(_197_),
    .A2(_198_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _457_ (.A1(\Datapath.k[12] ),
    .A2(net18),
    .B1(_082_),
    .B2(net4),
    .C1(_115_),
    .C2(\Datapath.k[13] ),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _458_ (.A1(_159_),
    .A2(_199_),
    .B(_200_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _459_ (.A1(\Datapath.k[13] ),
    .A2(\Datapath.k[12] ),
    .Z(_201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _460_ (.A1(\Datapath.k[12] ),
    .A2(\Datapath.k[11] ),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _461_ (.A1(_197_),
    .A2(_198_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _462_ (.A1(_202_),
    .A2(_203_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _463_ (.A1(_201_),
    .A2(_204_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _464_ (.I0(\Datapath.k[14] ),
    .I1(net5),
    .I2(_205_),
    .I3(\Datapath.k[13] ),
    .S0(_080_),
    .S1(_059_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _465_ (.I(_206_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _466_ (.A1(\Datapath.k[14] ),
    .A2(\Datapath.k[13] ),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _467_ (.A1(_197_),
    .A2(_198_),
    .A3(_201_),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _468_ (.A1(\Datapath.k[13] ),
    .A2(\Datapath.k[11] ),
    .B(\Datapath.k[12] ),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _469_ (.A1(_208_),
    .A2(_209_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _470_ (.A1(_207_),
    .A2(_210_),
    .Z(_211_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _471_ (.I0(\Datapath.k[15] ),
    .I1(net6),
    .I2(_211_),
    .I3(\Datapath.k[14] ),
    .S0(_080_),
    .S1(_059_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _472_ (.I(_212_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _473_ (.A1(\Datapath.k[15] ),
    .A2(\Datapath.k[14] ),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _474_ (.I(_207_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _475_ (.A1(_208_),
    .A2(_209_),
    .B(_214_),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _476_ (.A1(\Datapath.k[14] ),
    .A2(\Datapath.k[13] ),
    .B(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _477_ (.A1(_213_),
    .A2(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _478_ (.I0(\Datapath.k[16] ),
    .I1(net7),
    .I2(_217_),
    .I3(\Datapath.k[15] ),
    .S0(_080_),
    .S1(_059_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _479_ (.I(_218_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _480_ (.A1(\Datapath.k[16] ),
    .A2(\Datapath.k[15] ),
    .Z(_219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _481_ (.A1(_207_),
    .A2(_213_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _482_ (.A1(_209_),
    .A2(_220_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _483_ (.A1(_198_),
    .A2(_201_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _484_ (.A1(_193_),
    .A2(_196_),
    .B(_222_),
    .C(_220_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _485_ (.A1(\Datapath.k[15] ),
    .A2(\Datapath.k[13] ),
    .B(\Datapath.k[14] ),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _486_ (.I(_224_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _487_ (.A1(_219_),
    .A2(_221_),
    .A3(_223_),
    .A4(_225_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _488_ (.A1(_221_),
    .A2(_223_),
    .A3(_225_),
    .B(_219_),
    .ZN(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _489_ (.A1(_159_),
    .A2(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _490_ (.A1(\Datapath.k[17] ),
    .A2(_036_),
    .B1(_037_),
    .B2(\Datapath.k[16] ),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _491_ (.A1(_226_),
    .A2(_228_),
    .B(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _492_ (.A1(_082_),
    .A2(_230_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _493_ (.I(_231_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _494_ (.A1(\Datapath.k[18] ),
    .A2(_055_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _495_ (.A1(\Datapath.k[17] ),
    .A2(_055_),
    .B(_059_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _496_ (.A1(\Datapath.k[16] ),
    .A2(\Datapath.k[15] ),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _497_ (.A1(_234_),
    .A2(_227_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _498_ (.A1(\Datapath.k[17] ),
    .A2(\Datapath.k[16] ),
    .A3(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _499_ (.A1(_232_),
    .A2(_233_),
    .B1(_236_),
    .B2(_159_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _500_ (.A1(\Datapath.k[17] ),
    .A2(\Datapath.k[16] ),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _501_ (.A1(_069_),
    .A2(_227_),
    .B(_237_),
    .C(_234_),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _502_ (.A1(\Datapath.k[18] ),
    .A2(\Datapath.k[17] ),
    .A3(_238_),
    .Z(_239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _503_ (.A1(\Datapath.k[19] ),
    .A2(_036_),
    .B1(_159_),
    .B2(_239_),
    .C1(_037_),
    .C2(\Datapath.k[18] ),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _504_ (.A1(_061_),
    .A2(_240_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _505_ (.A1(\Datapath.k[18] ),
    .A2(\Datapath.k[17] ),
    .Z(_241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _506_ (.A1(\Datapath.k[18] ),
    .A2(\Datapath.k[17] ),
    .Z(_242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _507_ (.A1(_241_),
    .A2(_238_),
    .B(_242_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _508_ (.A1(\Datapath.k[19] ),
    .A2(\Datapath.k[18] ),
    .A3(_243_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _509_ (.A1(\Datapath.k[19] ),
    .A2(_037_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _510_ (.A1(_128_),
    .A2(_244_),
    .B(_245_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _511_ (.D(_000_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _512_ (.D(_001_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _513_ (.D(_002_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _514_ (.D(_003_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _515_ (.D(_004_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _516_ (.D(_005_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _517_ (.D(_006_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _518_ (.D(_007_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _519_ (.D(_008_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _520_ (.D(_009_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _521_ (.D(_010_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _522_ (.D(_011_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _523_ (.D(_012_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.i[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _524_ (.D(_013_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _525_ (.D(_014_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _526_ (.D(_015_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.i[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _527_ (.D(_016_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _528_ (.D(_017_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _529_ (.D(_018_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _530_ (.D(_019_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _531_ (.D(_020_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _532_ (.D(_021_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _533_ (.D(_022_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _534_ (.D(_023_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _535_ (.D(_024_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _536_ (.D(_025_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\Datapath.k[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _537_ (.D(_026_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _538_ (.D(_027_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _539_ (.D(_028_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _540_ (.D(_029_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _541_ (.D(_030_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _542_ (.D(_031_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _543_ (.D(_032_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _544_ (.D(_033_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _545_ (.D(_034_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _546_ (.D(_035_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _547_ (.D(\FSM.NS[0] ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\FSM.CS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _548_ (.D(\FSM.NS[1] ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(co[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(co[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(co[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(co[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(co[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(co[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(co[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(co[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(co[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(co[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(co[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(co[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(co[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(co[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(co[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(co[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(st),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(bs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(x[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(x[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(x[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(x[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(x[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(x[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(x[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(x[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(x[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(x[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(x[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(x[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(x[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(x[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(x[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(x[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A3 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__A1 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A2 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__A1 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__A1 (.I(\Datapath.i[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__A1 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__A1 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A1 (.I(\Datapath.i[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A2 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A1 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A1 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__A1 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A1 (.I(\Datapath.i[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A1 (.I(\Datapath.i[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__B (.I(\Datapath.i[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__A1 (.I(\Datapath.i[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__A2 (.I(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__A1 (.I(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__A1 (.I(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__A1 (.I(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__A1 (.I(\Datapath.i[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__A1 (.I(\Datapath.i[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__B (.I(\Datapath.i[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(\Datapath.i[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__A1 (.I(\Datapath.i[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__A1 (.I(\Datapath.i[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A2 (.I(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__B2 (.I(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A1 (.I(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A1 (.I(\Datapath.i[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A1 (.I(\Datapath.i[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A1 (.I(\Datapath.i[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A1 (.I(\Datapath.i[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A1 (.I(\Datapath.i[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__A1 (.I(\Datapath.i[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__A1 (.I(\Datapath.i[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A3 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A1 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__A1 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A1 (.I(\Datapath.i[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A2 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A1 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A1 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__A1 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A1 (.I(\Datapath.i[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A1 (.I(\Datapath.i[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__B (.I(\Datapath.i[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A1 (.I(\Datapath.i[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A2 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A1 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__A1 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A1 (.I(\Datapath.i[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A1 (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A1 (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__A1 (.I(\Datapath.i[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A1 (.I(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__A1 (.I(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A1 (.I(\Datapath.i[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__I (.I(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A3 (.I(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__A2 (.I(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A1 (.I(\Datapath.k[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A2 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__A1 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A1 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__A2 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__I3 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A1 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A2 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A2 (.I(\Datapath.k[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A2 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A2 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A2 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__I0 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A1 (.I(\Datapath.k[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__B (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A1 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A2 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A1 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A1 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A2 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A2 (.I(\Datapath.k[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A2 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__A2 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A1 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A2 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I3 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A1 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__C2 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A1 (.I(\Datapath.k[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__B (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__A1 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A2 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I3 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A1 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I0 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A4 (.I(\Datapath.k[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__A2 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A1 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A2 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I3 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__A1 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I0 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A3 (.I(\Datapath.k[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__A2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__A1 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__B2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__A1 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I0 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(\Datapath.k[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A2 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__500__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__498__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A1 (.I(\Datapath.k[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A2 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__506__A1 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A1 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__C2 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A1 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A1 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A2 (.I(\Datapath.k[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A1 (.I(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A1 (.I(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A1 (.I(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A1 (.I(\Datapath.k[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A2 (.I(\Datapath.k[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__A2 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A2 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__A1 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__A1 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__A1 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__I (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A2 (.I(\Datapath.k[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__A2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__B2 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A1 (.I(\Datapath.k[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__I (.I(\Datapath.k[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A2 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A2 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A1 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__C2 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A3 (.I(\Datapath.k[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A1 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A2 (.I(\Datapath.k[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__A2 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A2 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__B2 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A1 (.I(\Datapath.k[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A2 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__A2 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__A1 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__A2 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__A2 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A4 (.I(\Datapath.k[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__I (.I(\FSM.CS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A4 (.I(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__I (.I(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A2 (.I(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__I (.I(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A2 (.I(\FSM.CS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__547__D (.I(\FSM.NS[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__D (.I(\FSM.NS[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__D (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__D (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__D (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__D (.I(_003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__D (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__D (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__D (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__D (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__D (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__D (.I(_010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__D (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__D (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__D (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__D (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__D (.I(_015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__D (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__D (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__D (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__D (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__D (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__D (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__D (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__D (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__D (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__D (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__D (.I(_031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__D (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__D (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__D (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__I (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A1 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__C1 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__B1 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__C (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__I (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__B (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__I (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__B (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__B (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__B (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__B (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A3 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__B2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__A1 (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A1 (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A1 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__I (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__B (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__S1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__S1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__S1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__S1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__409__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__B (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__374__S (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__B1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__B1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__B1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__B (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__B (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__B (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__I (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__B1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__B2 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__A2 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__B1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__B2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A1 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A4 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A2 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__C2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A3 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A2 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A1 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A1 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A3 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__395__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__388__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__374__I0 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A4 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A3 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A4 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__B1 (.I(_078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__I (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__S0 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__S0 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__S0 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__S0 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__A1 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__B2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A2 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__A1 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__492__A1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__B1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__B1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__B1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__B1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__A1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__B (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__B (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__B1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A4 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A2 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__A2 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A3 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A2 (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A2 (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__A2 (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__A1 (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__I (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A3 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__A2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__A3 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A2 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__A2 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A1 (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A2 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__A2 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__A2 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__A3 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__A2 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A3 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A2 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A2 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__A2 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__A3 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__B (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__I (.I(_103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__A3 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__A2 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__A2 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__A2 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__A3 (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__B (.I(_106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__A2 (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__A2 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__A3 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__A2 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__B1 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__A2 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__A1 (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__A1 (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__C1 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__C1 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__B1 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__C1 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__B1 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__A2 (.I(_115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__A2 (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__B1 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__B2 (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__B2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__A1 (.I(_128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__A1 (.I(_128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__383__A2 (.I(_133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__A1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__A2 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A2 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__A2 (.I(_139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__400__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__C (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A4 (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A1 (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A1 (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__A2 (.I(_154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__407__A2 (.I(_154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__B (.I(_155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__411__A1 (.I(_156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__B1 (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__499__B2 (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A1 (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A1 (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__A1 (.I(_159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A2 (.I(_174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__431__B (.I(_176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__I (.I(_183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A1 (.I(_193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A2 (.I(_199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__481__A1 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__I (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__A1 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__C (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A1 (.I(_234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__A2 (.I(_238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A3 (.I(_238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__B2 (.I(_239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__A2 (.I(_240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(co[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(co[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(co[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(co[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(co[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(co[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(co[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(co[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(co[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(co[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(co[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(co[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(co[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(co[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(co[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(co[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(st));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__I1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A3 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__B2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A4 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__471__I1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A3 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A4 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__B1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A3 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__375__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A4 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__B2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__392__B2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A3 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__B2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__A4 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__B2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__B2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__C (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__C (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__541__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__CLK (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__518__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__524__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__527__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__543__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__CLK (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__513__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__547__CLK (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__516__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__539__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__548__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_687 ();
endmodule

