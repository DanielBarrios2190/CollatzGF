* NGSPICE file created from collatz.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

.subckt collatz bs clk co[0] co[10] co[11] co[12] co[13] co[14] co[15] co[1] co[2]
+ co[3] co[4] co[5] co[6] co[7] co[8] co[9] st vdd vss x[0] x[10] x[11] x[12] x[13]
+ x[14] x[15] x[1] x[2] x[3] x[4] x[5] x[6] x[7] x[8] x[9]
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__338__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__510__A1 _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_501_ _069_ _227_ _237_ _234_ _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_432_ Datapath.k\[10\] _070_ _177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_294_ net15 net16 net2 net3 _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_363_ _114_ _115_ _116_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__329__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__501__A1 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_346_ Datapath.i\[12\] Datapath.i\[11\] _101_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_415_ _144_ _145_ _143_ _152_ _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_277_ _052_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__410__B1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__401__B1 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__529__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_329_ _061_ _092_ _093_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__464__I0 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__392__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__383__A2 _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__365__A2 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 net20 x[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 x[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__292__A1 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__283__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__360__I Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_500_ Datapath.k\[17\] Datapath.k\[16\] _237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__274__A1 Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_362_ _059_ Datapath.k\[1\] net8 _061_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_431_ _169_ _175_ _176_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_293_ _062_ net8 net9 net10 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__501__A2 _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__256__A1 Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__495__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__247__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_345_ Datapath.i\[11\] _101_ Datapath.i\[12\] _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_414_ _072_ _131_ _160_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_276_ Datapath.i\[13\] _039_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__410__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__410__B2 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__401__B2 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__401__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__468__A1 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_328_ Datapath.i\[6\] Datapath.i\[5\] Datapath.i\[4\] _087_ _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_259_ _043_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__459__A1 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__464__I1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__519__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__359__B1 _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I co[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 x[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 x[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__292__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__347__A3 _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I co[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__283__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__338__A3 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__274__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_292_ net11 net12 net13 net14 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_430_ _070_ _037_ _060_ net16 _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_361_ _036_ _055_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__329__A3 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__256__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__281__I _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__495__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__247__A2 FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_413_ _129_ _136_ _143_ _152_ _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_344_ _103_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_275_ _051_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__410__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__401__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__468__A2 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_327_ Datapath.i\[5\] _088_ Datapath.i\[6\] _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_258_ Datapath.i\[4\] _039_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__459__A2 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__395__A1 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__386__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__310__A1 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__377__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__368__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__359__B2 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__359__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput22 net22 x[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 x[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__292__A3 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__408__B _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__504__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__369__I Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__279__I _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_291_ _057_ _063_ FSM.NS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_360_ Datapath.k\[2\] _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_489_ _159_ _227_ _228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_412_ _036_ _080_ _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_343_ Datapath.i\[11\] _101_ _102_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_274_ Datapath.i\[12\] _039_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_326_ _091_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_257_ _042_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__395__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__386__A2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__542__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__310__A2 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__464__I3 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_309_ FSM.CS\[1\] _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__377__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__368__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__359__A2 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__295__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput23 net23 x[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 x[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__292__A4 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__504__A2 _240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__268__A1 Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__440__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__334__B _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_290_ _059_ net17 _061_ _062_ _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__498__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__422__A1 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_488_ _221_ _223_ _225_ _219_ _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__489__A1 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_411_ _156_ _157_ _158_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_342_ Datapath.i\[11\] _101_ _060_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__404__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_273_ _050_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_325_ Datapath.i\[5\] _088_ _090_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__313__B1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_256_ Datapath.i\[3\] _039_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__342__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_308_ _079_ FSM.NS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__295__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__532__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput24 net24 x[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__268__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__440__A2 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__498__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_487_ _219_ _221_ _223_ _225_ _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__489__A2 _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I co[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__413__A2 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__345__B Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__511__D _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__404__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_341_ _061_ _100_ _101_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_410_ Datapath.k\[7\] _037_ _060_ net14 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_272_ Datapath.i\[11\] _039_ _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__340__A1 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_539_ _028_ clknet_2_3__leaf_clk Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__331__A1 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__398__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__322__A1 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__389__A1 _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_324_ Datapath.i\[5\] _088_ _060_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_255_ _041_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__313__B2 Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__313__A1 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__304__A1 Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_307_ _061_ _068_ _078_ _055_ _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__295__A3 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__348__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__514__D _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 x[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_486_ _224_ _225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__522__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_340_ Datapath.i\[10\] _099_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__545__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_271_ _049_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__340__A2 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_538_ _027_ clknet_2_1__leaf_clk Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__446__B _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_469_ _208_ _209_ _210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__331__A2 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__398__A2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__522__D _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__322__A2 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_323_ _088_ _089_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_254_ Datapath.i\[2\] _039_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__313__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__304__A2 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__517__D _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_306_ _069_ _071_ _075_ _077_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__470__A1 _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__295__A4 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__507__A2 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__530__D _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 x[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__434__A1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__416__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__525__D _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__407__A1 _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_485_ Datapath.k\[15\] Datapath.k\[13\] Datapath.k\[14\] _224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__413__A4 _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_270_ Datapath.i\[10\] _039_ _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_468_ Datapath.k\[13\] Datapath.k\[11\] Datapath.k\[12\] _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_537_ _026_ clknet_2_0__leaf_clk Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_399_ _143_ _147_ _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__478__S0 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__307__B1 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__512__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_322_ Datapath.i\[4\] _087_ _082_ _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_253_ _040_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__301__I Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__304__A3 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__535__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__533__D _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_305_ Datapath.k\[0\] _056_ _076_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__528__D _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 x[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__434__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__370__A1 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__361__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__416__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__352__A1 Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__541__D _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__407__A2 _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_484_ _193_ _196_ _222_ _220_ _223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__343__A1 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__334__A1 Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__325__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_467_ _197_ _198_ _201_ _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_536_ _025_ clknet_2_2__leaf_clk Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_398_ Datapath.k\[5\] _073_ _137_ _146_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__316__A1 Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__478__S1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__307__B2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__307__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_321_ Datapath.i\[4\] _087_ _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_252_ Datapath.i\[1\] _039_ _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_519_ _008_ clknet_2_0__leaf_clk Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__304__A4 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_304_ Datapath.k\[19\] Datapath.k\[18\] Datapath.k\[15\] Datapath.k\[14\] _076_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__468__B Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__544__D _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__525__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 x[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__548__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__370__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__361__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__375__C _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__391__B _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__352__A2 Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_483_ _198_ _201_ _222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__343__A2 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__270__A1 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__325__A2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_535_ _024_ clknet_2_3__leaf_clk Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_466_ Datapath.k\[14\] Datapath.k\[13\] _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_397_ _144_ _145_ _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__316__A2 Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__252__A1 Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__307__A2 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__547__D FSM.NS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_320_ _061_ _086_ _087_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_251_ _037_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_518_ _007_ clknet_2_1__leaf_clk Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_449_ _166_ _170_ _177_ _184_ _192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__473__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_303_ Datapath.k\[7\] Datapath.k\[6\] _072_ _074_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__455__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__446__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput18 net18 bs vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net29 x[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__419__A1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__352__A3 _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__515__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_482_ _209_ _220_ _221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__538__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__270__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_465_ _206_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_534_ _023_ clknet_2_2__leaf_clk Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_396_ Datapath.k\[5\] _073_ _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__316__A3 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__252__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_250_ _038_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_517_ _006_ clknet_2_0__leaf_clk Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_448_ _189_ _190_ _191_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__326__I _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_379_ Datapath.k\[3\] Datapath.k\[2\] _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__473__A2 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_302_ Datapath.k\[11\] Datapath.k\[10\] Datapath.k\[5\] _073_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__455__A2 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__391__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__446__A2 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__373__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__495__B _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__364__A1 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 x[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__419__A2 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__355__A1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__346__A1 Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__337__A1 Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_481_ _207_ _213_ _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__328__A1 Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__500__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__319__A1 Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_464_ Datapath.k\[14\] net5 _205_ Datapath.k\[13\] _080_ _059_ _206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_533_ _022_ clknet_2_2__leaf_clk Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__316__A4 FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_395_ _073_ Datapath.k\[3\] _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_516_ _005_ clknet_2_3__leaf_clk Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__528__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_447_ Datapath.k\[11\] _037_ _060_ net3 _191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_378_ _073_ Datapath.k\[3\] _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_73_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_301_ Datapath.k\[4\] _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__391__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__373__A2 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__364__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I co[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__355__A2 _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__291__A1 _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__346__A2 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__503__C1 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input8_I co[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__337__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_480_ Datapath.k\[16\] Datapath.k\[15\] _219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__328__A2 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__264__A1 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__494__A1 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_463_ _201_ _204_ _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_532_ _021_ clknet_2_0__leaf_clk Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_394_ Datapath.k\[6\] Datapath.k\[5\] _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__485__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__476__A1 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__400__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_515_ _004_ clknet_2_3__leaf_clk Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_377_ _059_ _055_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_446_ _059_ Datapath.k\[12\] _055_ _190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__458__A1 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_300_ Datapath.k\[3\] Datapath.k\[2\] _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__471__S0 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_429_ _036_ _174_ _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput1 co[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__367__B1 _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__374__S _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__364__A3 Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__503__B1 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__346__A3 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__503__C2 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__328__A3 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__264__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__421__C1 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__310__B _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__494__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_531_ _020_ clknet_2_3__leaf_clk Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_462_ _202_ _203_ _204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_393_ _140_ _141_ _142_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__485__A2 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__476__A2 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__400__A2 _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_514_ _003_ clknet_2_3__leaf_clk Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_376_ _120_ _127_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_445_ _036_ _188_ _189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__458__A2 _199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__394__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__385__A1 _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_428_ _170_ _173_ _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__471__S1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_359_ _062_ _061_ _112_ _080_ _113_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__300__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput2 co[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__367__A1 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__367__B2 _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__358__A1 _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__349__A1 Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__503__A1 Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__503__B2 _239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__430__B1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__328__A4 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__421__B1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__421__C2 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_530_ _019_ clknet_2_3__leaf_clk Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_461_ _197_ _198_ _203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_392_ Datapath.k\[5\] _037_ _061_ net12 _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__282__I FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_513_ _002_ clknet_2_2__leaf_clk Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_444_ _184_ _187_ _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_375_ _080_ net10 _082_ _126_ _037_ _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__394__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__385__A2 _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_427_ _165_ _171_ _172_ _173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_358_ _057_ _112_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__541__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_289_ net1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__300__A2 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 co[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__358__A2 _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__294__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__349__A2 _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__276__A1 Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__503__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__324__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__258__A1 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input14_I co[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__430__A1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__430__B2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__285__I _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__497__A1 _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__249__A1 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__421__A1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__421__B2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__409__B _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I co[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__412__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__501__C _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_460_ Datapath.k\[12\] Datapath.k\[11\] _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_391_ _059_ Datapath.k\[6\] _055_ _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_512_ _001_ clknet_2_2__leaf_clk Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_443_ _185_ _181_ _186_ _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_374_ _073_ _125_ _059_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_426_ Datapath.k\[8\] Datapath.k\[7\] _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_357_ _036_ Datapath.k\[0\] _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_288_ _060_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 co[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__327__B Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__288__I _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__438__S0 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__294__A2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_409_ _059_ Datapath.k\[8\] _055_ _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__531__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__276__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__258__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__430__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__497__A2 _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__249__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__421__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__412__A2 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_390_ _036_ _139_ _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__330__A1 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__321__A1 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_511_ _000_ clknet_2_3__leaf_clk Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_373_ Datapath.k\[3\] Datapath.k\[2\] _124_ _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_442_ Datapath.k\[10\] _070_ _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__388__A1 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__312__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__379__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__303__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_287_ _058_ FSM.CS\[1\] _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_356_ _111_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_425_ _166_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput5 co[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__343__B _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__438__S1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__294__A3 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ _152_ _154_ _155_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_339_ Datapath.i\[10\] _099_ _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__506__A1 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__521__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__351__B Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__478__I0 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__544__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__330__A2 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__512__D _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__321__A2 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_510_ _128_ _244_ _245_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_441_ Datapath.k\[10\] _070_ _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__388__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_372_ _121_ _122_ _123_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__312__A2 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__379__A2 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__303__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_424_ _070_ Datapath.k\[8\] _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_355_ _082_ _110_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_286_ _058_ _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__297__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 co[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__460__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__294__A4 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__451__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_338_ _061_ _098_ _099_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_407_ _152_ _154_ _059_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__506__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_269_ _048_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__442__A1 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__520__D _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__424__A1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__349__B _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__515__D _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I co[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__478__I1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I co[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_371_ Datapath.k\[2\] Datapath.k\[1\] _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_440_ Datapath.k\[11\] Datapath.k\[10\] _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__511__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__303__A3 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__523__D _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__534__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_423_ _059_ Datapath.k\[10\] _055_ _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_354_ Datapath.i\[15\] _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_285_ _036_ _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__297__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 co[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__460__A2 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__518__D _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__451__A2 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_337_ Datapath.i\[9\] _096_ _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_406_ _143_ _147_ _153_ _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_268_ Datapath.i\[9\] _039_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__442__A2 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__424__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput10 co[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__531__D _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__351__A1 Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__342__A1 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__333__A1 Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__526__D _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__324__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__315__A1 Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__306__A1 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__490__B1 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_370_ Datapath.k\[2\] Datapath.k\[1\] _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_499_ _232_ _233_ _236_ _159_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_422_ _159_ _167_ _168_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_353_ _061_ _108_ _109_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_284_ _055_ _056_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 co[1] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__509__A1 Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_336_ Datapath.i\[9\] _096_ _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_405_ Datapath.k\[6\] Datapath.k\[5\] _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_267_ _047_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__524__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__547__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput11 co[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_319_ Datapath.i\[3\] _085_ _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__351__A2 _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__342__A2 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__333__A2 Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__542__D _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__478__I3 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__324__A2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__260__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__315__A2 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__306__A2 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__490__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__490__B2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__537__D _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__481__A1 _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_498_ Datapath.k\[17\] Datapath.k\[16\] _235_ _236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_421_ Datapath.k\[8\] net18 _082_ net15 _115_ _070_ _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_85_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_352_ Datapath.i\[14\] Datapath.i\[13\] _105_ _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_81_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_283_ _036_ Datapath.k\[1\] _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 co[2] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__454__A1 _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__509__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__445__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__436__A1 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_404_ Datapath.k\[7\] Datapath.k\[6\] _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_335_ _096_ _097_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_266_ Datapath.i\[8\] _039_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__409__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__308__I _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 co[5] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_318_ Datapath.i\[3\] _085_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_249_ Datapath.i\[0\] _037_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__514__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__333__A3 _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__537__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__260__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__306__A3 _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I co[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__490__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_497_ _234_ _227_ _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__457__C1 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I co[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__548__D FSM.NS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_351_ Datapath.i\[13\] _105_ Datapath.i\[14\] _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_420_ _165_ _166_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_282_ FSM.CS\[1\] _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__390__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__381__A1 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__436__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_334_ Datapath.i\[8\] _095_ _082_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_403_ _149_ _150_ _151_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_265_ _046_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__485__B Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__363__A1 _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__354__A1 Datapath.i\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__409__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__290__B1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 co[6] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_317_ _061_ _084_ _085_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__345__A1 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_248_ _037_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_84_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__336__A1 Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__327__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__318__A1 Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__306__A4 _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_496_ Datapath.k\[16\] Datapath.k\[15\] _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__457__C2 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__457__B1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__527__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__471__I0 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_350_ _107_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__384__C1 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_281_ _054_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_548_ FSM.NS\[1\] clknet_2_3__leaf_clk FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_479_ _218_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__390__A2 _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__381__A2 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_333_ Datapath.i\[8\] Datapath.i\[7\] _093_ _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_402_ Datapath.k\[6\] _037_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_264_ Datapath.i\[7\] _039_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__363__A2 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__354__A2 _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__290__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__290__B2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput14 co[7] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_316_ Datapath.i\[2\] Datapath.i\[1\] Datapath.i\[0\] FSM.CS\[1\] _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_247_ _036_ FSM.CS\[1\] _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__345__A2 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__336__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__250__I _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__272__A1 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__327__A2 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__254__A1 Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__484__A1 _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__466__A1 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_495_ Datapath.k\[17\] _055_ _059_ _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__457__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__457__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__471__I1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_280_ Datapath.i\[15\] _037_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__384__B1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__384__C2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_547_ FSM.NS\[0\] clknet_2_2__leaf_clk FSM.CS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_478_ Datapath.k\[16\] net7 _217_ Datapath.k\[15\] _080_ _059_ _218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__375__B1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__366__B1 _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_401_ _055_ net13 _115_ Datapath.k\[7\] net18 _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_76_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_332_ _061_ _094_ _095_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_263_ _045_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__517__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__248__I _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__290__A2 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput15 co[8] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_315_ Datapath.i\[2\] _081_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_246_ FSM.CS\[0\] _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__272__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__254__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__466__A2 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_494_ Datapath.k\[18\] _055_ _232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__457__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__384__B2 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__384__A1 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_546_ _035_ clknet_2_0__leaf_clk Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_477_ _213_ _216_ _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__375__A1 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__375__B2 _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__366__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__366__B2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_331_ Datapath.i\[7\] _093_ _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_400_ _036_ _148_ _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__357__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_262_ Datapath.i\[6\] _039_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_529_ _018_ clknet_2_0__leaf_clk Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__348__A1 Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__339__A1 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__439__I _183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_314_ _081_ _083_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 co[9] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__502__A1 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_493_ _231_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__471__I3 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__384__A2 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_545_ _034_ clknet_2_1__leaf_clk Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_476_ Datapath.k\[14\] Datapath.k\[13\] _215_ _216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__375__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__438__I0 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__540__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__366__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_330_ Datapath.i\[7\] _093_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__357__A2 Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_261_ _044_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__293__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_459_ Datapath.k\[13\] Datapath.k\[12\] _201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_528_ _017_ clknet_2_2__leaf_clk Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__348__A2 _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__284__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__339__A2 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_313_ Datapath.i\[0\] _055_ _082_ Datapath.i\[1\] _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 st net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__502__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__266__A1 Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__496__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__411__A1 _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__402__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__401__C net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_492_ _082_ _230_ _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__322__B _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__464__S0 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_544_ _033_ clknet_2_3__leaf_clk Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_475_ _208_ _209_ _214_ _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__407__B _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__438__I1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__374__I0 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_260_ Datapath.i\[5\] _039_ _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__293__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_527_ _016_ clknet_2_1__leaf_clk Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_458_ _159_ _199_ _200_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_389_ _136_ _138_ _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__284__A2 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_312_ _036_ _080_ _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__502__A3 _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__530__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__266__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__496__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__402__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__286__I _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__396__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__320__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_491_ _226_ _228_ _229_ _230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__311__A1 Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__378__A1 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__302__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__464__S1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_543_ _032_ clknet_2_1__leaf_clk Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__474__I _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_474_ _207_ _214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__423__B _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__293__A3 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_526_ _015_ clknet_2_2__leaf_clk Datapath.i\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_457_ Datapath.k\[12\] net18 _082_ net4 _115_ Datapath.k\[13\] _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_82_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_388_ _073_ Datapath.k\[3\] _137_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__505__A1 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__289__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_311_ Datapath.i\[1\] Datapath.i\[0\] _055_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_509_ Datapath.k\[19\] _037_ _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__415__C _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__431__B _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input17_I st vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__520__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I co[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__396__A2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__543__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_490_ Datapath.k\[17\] _036_ _037_ Datapath.k\[16\] _229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__311__A2 Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__378__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__302__A2 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_542_ _031_ clknet_2_3__leaf_clk Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_473_ Datapath.k\[15\] Datapath.k\[14\] _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__296__A1 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__438__I3 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__287__A1 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__278__A1 Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__293__A4 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_456_ _197_ _198_ _199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_525_ _014_ clknet_2_2__leaf_clk Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_387_ _129_ _132_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__505__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__441__A1 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_310_ Datapath.i\[0\] _080_ _038_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__432__A1 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__499__B2 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__423__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_439_ _183_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_508_ Datapath.k\[19\] Datapath.k\[18\] _243_ _244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__414__A1 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__405__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__320__A3 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__311__A3 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__302__A3 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__513__D _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_472_ _212_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_541_ _030_ clknet_2_0__leaf_clk Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__533__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__287__A2 FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__278__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_524_ _013_ clknet_2_1__leaf_clk Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_455_ Datapath.k\[12\] Datapath.k\[11\] _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_386_ Datapath.k\[5\] _073_ _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_72_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__441__A2 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__432__A2 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__423__A2 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_438_ Datapath.k\[11\] net2 _182_ Datapath.k\[10\] _080_ _059_ _183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_507_ _241_ _238_ _242_ _243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_369_ Datapath.k\[0\] _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__414__A2 _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__521__D _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__405__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__341__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__332__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__516__D _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__323__A1 _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__314__A1 _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__305__A1 Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__A4 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_540_ _029_ clknet_2_1__leaf_clk Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_471_ Datapath.k\[15\] net6 _211_ Datapath.k\[14\] _080_ _059_ _212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__508__A1 Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__524__D _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_523_ _012_ clknet_2_3__leaf_clk Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_454_ _193_ _196_ _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_385_ _134_ _135_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__523__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_506_ Datapath.k\[18\] Datapath.k\[17\] _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_368_ Datapath.k\[3\] net18 _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_437_ _177_ _181_ _182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_299_ Datapath.k\[13\] Datapath.k\[12\] _070_ Datapath.k\[8\] _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__546__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__341__A2 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__532__D _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__305__A2 _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input15_I co[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__527__D _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__480__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__299__A1 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I co[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_470_ _207_ _210_ _211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__296__A4 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__508__A2 Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__540__D _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_522_ _011_ clknet_2_1__leaf_clk Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_453_ _186_ _194_ _195_ _196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_384_ _073_ net18 _082_ net11 _115_ Datapath.k\[5\] _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_41_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__426__A1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__B1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__408__A1 _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_436_ _070_ Datapath.k\[8\] _178_ _180_ _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_505_ Datapath.k\[18\] Datapath.k\[17\] _241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_298_ Datapath.k\[9\] _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_367_ _114_ net18 _118_ _119_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__341__A3 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_419_ Datapath.k\[8\] Datapath.k\[7\] _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__513__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__366__C net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__536__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__543__D _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__480__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__299__A2 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__538__D _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_383_ _128_ _133_ _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_521_ _010_ clknet_2_3__leaf_clk Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_452_ _177_ _180_ _184_ _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__371__A1 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__426__A2 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__362__A1 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__362__B2 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__353__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__408__A2 _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_504_ _061_ _240_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_366_ _055_ net9 _115_ Datapath.k\[3\] net18 _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_435_ _172_ _179_ _180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_297_ Datapath.k\[17\] Datapath.k\[16\] _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__335__A1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__546__D _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__309__I FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_349_ Datapath.i\[13\] _105_ _106_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_418_ _161_ _162_ _164_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__317__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__299__A3 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__447__B1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__526__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_520_ _009_ clknet_2_1__leaf_clk Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_451_ Datapath.k\[11\] Datapath.k\[10\] _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_382_ _129_ _132_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__371__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__362__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__353__A2 _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_503_ Datapath.k\[19\] _036_ _159_ _239_ _037_ Datapath.k\[18\] _240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_296_ _064_ _065_ _066_ _067_ _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_434_ _070_ Datapath.k\[8\] _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_365_ _036_ _117_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__280__A1 Datapath.i\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__335__A2 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__262__A1 Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_417_ _153_ _163_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_348_ Datapath.i\[13\] _105_ _060_ _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_279_ _053_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__492__A1 _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__299__A4 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__392__B1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__447__B2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__447__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I co[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I co[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__429__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_450_ _161_ _162_ _164_ _192_ _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_381_ _072_ _131_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__516__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__353__A3 _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_502_ Datapath.k\[18\] Datapath.k\[17\] _238_ _239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_433_ _165_ _171_ _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_295_ net4 net5 net6 net7 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_364_ Datapath.k\[2\] Datapath.k\[1\] Datapath.k\[0\] _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__539__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__280__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_416_ Datapath.k\[7\] Datapath.k\[6\] _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__262__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_347_ _061_ _104_ _105_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_278_ Datapath.i\[14\] _039_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__251__I _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__246__I FSM.CS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__392__B2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__392__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__447__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__383__A1 _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__429__A2 _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__365__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_380_ _121_ _122_ _130_ _123_ _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput30 net30 x[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__344__I _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__347__A1 _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

