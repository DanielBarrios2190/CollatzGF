* NGSPICE file created from collatz.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

.subckt collatz bs clk co[0] co[10] co[11] co[12] co[13] co[14] co[15] co[1] co[2]
+ co[3] co[4] co[5] co[6] co[7] co[8] co[9] st vdd vss x[0] x[10] x[11] x[12] x[13]
+ x[14] x[15] x[1] x[2] x[3] x[4] x[5] x[6] x[7] x[8] x[9]
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__510__A1 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__429__I _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_501_ _042_ _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_432_ _040_ _037_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_363_ _047_ Datapath.i\[5\] _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__568__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__559__A1 _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_415_ Datapath.k\[14\] _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_346_ _037_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_680_ _315_ _311_ _320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__717__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_732_ _025_ clknet_2_1__leaf_clk Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_594_ _080_ _075_ _241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_663_ _222_ _303_ _304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__677__A3 _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput20 net20 x[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 x[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_715_ _008_ clknet_2_3__leaf_clk Datapath.i\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__347__A2 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__595__A2 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__625__I _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_646_ Datapath.k\[15\] _103_ _038_ net6 _046_ _289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_577_ _222_ _225_ _226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__360__I _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_500_ _103_ Datapath.k\[1\] _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_362_ _048_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_431_ _074_ _104_ FSM.NS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_629_ _270_ _272_ _273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_345_ FSM.CS\[1\] _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_414_ Datapath.k\[15\] _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__477__A1 _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__640__A1 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__459__A1 _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__698__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__698__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__699__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__689__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_731_ _024_ clknet_2_1__leaf_clk Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_662_ _302_ _238_ _255_ _303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_593_ _221_ _238_ _239_ _240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input11_I co[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__589__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput21 net21 x[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 x[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_645_ _286_ _064_ _287_ _288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_714_ _007_ clknet_2_3__leaf_clk Datapath.i\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_576_ _223_ _224_ _225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__504__B1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I co[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__707__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__510__A3 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_361_ _047_ Datapath.i\[4\] _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_430_ _092_ _101_ _103_ _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_628_ _100_ _271_ _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_559_ _094_ _205_ _209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_413_ Datapath.k\[5\] Datapath.k\[4\] _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_344_ FSM.CS\[0\] _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__477__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__640__A2 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__631__A2 _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__395__A1 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__622__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__386__A1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__689__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__740__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__604__A2 _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__368__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__540__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_661_ _301_ _302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_592_ _224_ _232_ _239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_730_ _023_ clknet_2_1__leaf_clk Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__522__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__589__A1 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__513__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput22 net22 x[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 x[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_713_ _006_ clknet_2_2__leaf_clk Datapath.i\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_644_ _278_ _280_ _284_ _287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_575_ Datapath.k\[8\] Datapath.k\[7\] _224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__504__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__504__B2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_360_ _046_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_627_ Datapath.k\[13\] Datapath.k\[12\] _271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_558_ _204_ _207_ _208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_489_ _141_ Datapath.i\[13\] Datapath.i\[12\] Datapath.i\[11\] _149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__652__I _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_412_ Datapath.k\[0\] _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__631__A3 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__395__A2 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__386__A2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__368__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_660_ _277_ _300_ _301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_591_ _225_ _233_ _238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__390__I Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__522__A2 _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__589__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__513__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 x[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 x[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__730__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_712_ _005_ clknet_2_3__leaf_clk Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_643_ _281_ _285_ _286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_574_ _076_ _213_ _223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__504__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__431__A1 _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__498__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__670__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_488_ _056_ _145_ _148_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_626_ _261_ _262_ _269_ _270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_557_ _206_ _093_ _207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__489__A1 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__413__A1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_411_ _077_ _078_ _081_ _084_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_609_ _253_ _254_ _079_ _047_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__634__A1 _265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_590_ _236_ _237_ _075_ _158_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 x[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_642_ _284_ _285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_711_ _004_ clknet_2_3__leaf_clk Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_573_ _221_ _222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__431__A2 _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__670__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_625_ _263_ _269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_487_ _147_ _062_ _148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_556_ _205_ _206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I co[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__413__A2 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__720__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_410_ _082_ _083_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__743__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_608_ Datapath.k\[12\] _103_ _038_ net3 _046_ _254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_539_ net12 _120_ Datapath.k\[6\] _102_ _042_ _191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__634__A2 _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__543__A1 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__525__A1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__516__A1 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__507__A1 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__530__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 x[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_710_ _003_ clknet_2_2__leaf_clk Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_641_ _282_ _283_ _284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_572_ _217_ _220_ _221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_624_ _267_ _268_ _099_ _047_ _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_555_ Datapath.k\[7\] Datapath.k\[6\] _205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_486_ _146_ _147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__646__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_607_ _251_ _252_ _253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_538_ _185_ _188_ _189_ _190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_469_ _131_ _053_ _062_ _133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__398__A2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__561__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__710__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__623__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__733__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__470__A1 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__525__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__516__A2 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__507__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__443__A1 _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 x[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_640_ Datapath.k\[14\] Datapath.k\[13\] _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_571_ _218_ _192_ _219_ _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__407__A1 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_485_ _143_ _056_ _146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_623_ Datapath.k\[13\] _103_ _038_ net4 _046_ _268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_554_ _200_ _195_ _204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__646__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__489__A4 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__628__A1 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_537_ _185_ _188_ _060_ _189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_468_ _052_ _129_ _132_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_606_ _244_ _242_ _249_ _252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_399_ _060_ _037_ _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__398__A3 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__519__B1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__443__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__691__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__723__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 x[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__539__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_570_ _195_ _205_ _219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__370__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_699_ _336_ _337_ _121_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__361__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__416__A2 _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__407__A2 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_622_ _264_ _064_ _266_ _267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_484_ _141_ Datapath.i\[11\] _145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_553_ _201_ _202_ _203_ _158_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__646__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__582__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__628__A2 _271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_605_ _250_ _036_ _251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__564__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_398_ _070_ _060_ net1 _071_ _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_467_ _131_ _062_ _132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_536_ _187_ _087_ _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__619__A2 _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__555__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__546__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__537__A1 _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_519_ net10 _121_ Datapath.k\[4\] _102_ _042_ _173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__528__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__402__I Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__519__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__600__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput28 net28 x[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_698_ _042_ Datapath.k\[18\] Datapath.k\[19\] _060_ _337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__361__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__391__B _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__655__A3 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_621_ _260_ _265_ _266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_483_ _055_ _140_ _144_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_552_ Datapath.k\[6\] _203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__713__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__736__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__405__I Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_535_ _186_ _184_ _187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_604_ _244_ _242_ _249_ _250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_397_ net8 net9 net10 net11 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_466_ _128_ Datapath.i\[8\] Datapath.i\[7\] _131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__619__A3 _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__555__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__546__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_518_ _169_ _064_ _171_ _172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__537__A2 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_449_ _117_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__528__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__519__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__446__A1 _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__437__A1 _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__437__B2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__479__B _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__600__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput18 net18 bs vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net29 x[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__419__A1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__408__I Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_697_ _334_ _317_ _335_ _336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__656__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_551_ net13 _120_ Datapath.k\[7\] _102_ _046_ _202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_620_ _262_ _263_ _265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_482_ _143_ _062_ _144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__421__I Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_465_ _051_ _127_ _130_ _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_534_ Datapath.k\[5\] _186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_603_ _081_ _248_ _249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_396_ _069_ net5 net6 net7 _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_4_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__491__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__482__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_448_ _115_ Datapath.i\[4\] _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_517_ _165_ _162_ _170_ _171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_379_ Datapath.i\[13\] _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__726__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__464__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__455__A2 _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__391__A1 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__382__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__437__A2 _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__685__A2 _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__373__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__600__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 x[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__419__A2 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__424__I Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__355__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__594__A1 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_696_ _329_ _333_ _335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_481_ _142_ Datapath.i\[11\] Datapath.i\[10\] _143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_550_ _199_ _200_ _036_ _201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__500__A1 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_679_ _318_ _319_ _121_ _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_602_ Datapath.k\[11\] Datapath.k\[10\] _248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_464_ _129_ _062_ _130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_533_ _181_ _176_ _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_395_ _067_ _068_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_447_ _115_ Datapath.i\[4\] _062_ _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_378_ net18 _056_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_516_ _097_ _168_ _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__498__B _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__391__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__382__A2 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__373__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__716__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I co[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__355__A2 Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__739__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__440__I _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_695_ _329_ _333_ _334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_15_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I co[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_480_ _131_ _053_ _142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__500__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_678_ _047_ Datapath.k\[16\] Datapath.k\[17\] _060_ _319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_601_ _246_ _247_ _080_ _158_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_394_ net12 net13 net14 net15 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_532_ _182_ _183_ _184_ _158_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_463_ _128_ Datapath.i\[7\] _129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__703__A2 _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_515_ _167_ _097_ _168_ _169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_446_ _113_ _114_ _115_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_377_ Datapath.i\[12\] _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__630__A1 _270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__689__B Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__621__A1 _260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__612__A1 _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_429_ _102_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_5_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 co[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_3_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__438__I Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__530__B1 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__348__I _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__512__B1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_694_ _332_ _333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_677_ _313_ _315_ _317_ _318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__729__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_600_ Datapath.k\[11\] _103_ _038_ net2 _046_ _247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_531_ Datapath.k\[4\] _184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_17_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_393_ net16 net2 net3 net4 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_462_ _126_ _128_ _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_729_ _022_ clknet_2_1__leaf_clk Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__356__I _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__400__A2 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__467__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_514_ Datapath.k\[3\] Datapath.k\[2\] _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_445_ _113_ _045_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_376_ net18 _055_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__458__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__394__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__630__A2 _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__697__A2 _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__621__A2 _265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_428_ _073_ _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__376__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__612__A2 _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_359_ _041_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__603__A2 _248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 co[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_3_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__530__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__521__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__512__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_693_ _330_ _331_ _332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__503__A1 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_676_ _316_ _317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__552__I Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__494__A3 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_530_ net11 _120_ Datapath.k\[5\] _102_ _042_ _183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_461_ _127_ _128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_392_ net1 _062_ _063_ _066_ FSM.NS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__637__I _279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_659_ _284_ _293_ _300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_728_ _021_ clknet_2_1__leaf_clk Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__633__B1 _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__400__A3 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__624__B1 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_513_ _165_ _162_ _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_444_ _062_ Datapath.i\[3\] _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_375_ Datapath.i\[11\] _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__719__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__458__A3 _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__394__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_427_ _065_ _094_ _097_ _100_ _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_358_ net18 _045_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__376__A2 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 co[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__358__A2 _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__521__A2 Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__512__A2 _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_692_ Datapath.k\[18\] Datapath.k\[17\] _331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__503__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__375__I Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input14_I co[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_744_ FSM.NS\[1\] clknet_2_0__leaf_clk FSM.CS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_675_ _036_ _037_ _316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input6_I co[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__651__A1 _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_391_ _064_ _065_ _037_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_460_ _125_ Datapath.i\[6\] _127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_727_ _020_ clknet_2_0__leaf_clk Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_658_ _297_ _298_ _299_ _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_589_ Datapath.k\[10\] _103_ _038_ net16 _046_ _237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__633__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__563__I Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__624__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_512_ _160_ _166_ _096_ _158_ _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_374_ _054_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_443_ _110_ _037_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__551__B1 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_426_ _098_ _099_ _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_357_ Datapath.i\[3\] _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput4 co[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__709__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_409_ Datapath.k\[16\] _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__504__C _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_691_ Datapath.k\[18\] Datapath.k\[17\] _330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__430__B _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_743_ FSM.NS\[0\] clknet_2_0__leaf_clk FSM.CS\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_674_ _304_ _308_ _314_ _315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__476__I _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__479__A2 _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_390_ Datapath.k\[1\] _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_657_ _039_ Datapath.k\[15\] _299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_726_ _019_ clknet_2_0__leaf_clk Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_588_ _231_ _234_ _235_ _236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__397__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__742__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_511_ _164_ _036_ _165_ _166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__388__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_442_ _112_ _044_ _109_ _106_ _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_373_ _047_ Datapath.i\[10\] _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_709_ _002_ clknet_2_2__leaf_clk Datapath.i\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__551__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__394__A4 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__551__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__606__A2 _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__533__A1 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__433__B _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_425_ Datapath.k\[12\] _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_356_ _044_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput5 co[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_32_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__515__A1 _167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_408_ Datapath.k\[17\] _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__506__A1 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__389__I _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_690_ _309_ _327_ _328_ _329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__497__A3 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_742_ _035_ clknet_2_3__leaf_clk Datapath.k\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_673_ _312_ _314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_725_ _018_ clknet_2_0__leaf_clk Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_656_ Datapath.k\[16\] _103_ _038_ net7 _042_ _298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_587_ _231_ _234_ _060_ _235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__609__B1 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_510_ _161_ Datapath.k\[0\] _162_ _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_441_ _111_ _037_ _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_372_ net18 _053_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_708_ _001_ clknet_2_2__leaf_clk Datapath.i\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_639_ _089_ _098_ _282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_424_ Datapath.k\[13\] _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__533__A2 _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_355_ _042_ Datapath.i\[2\] _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__732__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 co[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__608__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__460__A1 _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__515__A2 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_407_ _079_ _080_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__506__A2 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__442__B2 _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__433__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__681__A1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_741_ _034_ clknet_2_3__leaf_clk Datapath.k\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_672_ _309_ _312_ _313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__581__B1 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__636__A1 _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I co[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__627__A1 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_724_ _017_ clknet_2_0__leaf_clk Datapath.k\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_586_ _233_ _234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_655_ _295_ _296_ _064_ _297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__618__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I co[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__609__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__537__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_371_ Datapath.i\[9\] _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_440_ _110_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_707_ _000_ clknet_2_2__leaf_clk Datapath.i\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_638_ _278_ _280_ _281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_569_ _215_ _218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__447__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_423_ _095_ _096_ _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_354_ _043_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 co[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__515__A3 _168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__451__A2 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_406_ Datapath.k\[10\] _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_24_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__442__A2 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__681__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__433__A2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__722__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 co[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__654__A2 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_740_ _033_ clknet_2_3__leaf_clk Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_671_ _310_ _311_ _312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__590__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__645__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__581__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__632__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__581__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__636__A2 _271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__572__A1 _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__627__A2 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_723_ _016_ clknet_2_0__leaf_clk Datapath.k\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_654_ _286_ _283_ _293_ _296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_585_ _077_ _232_ _233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__618__A2 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_370_ net18 _052_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_637_ _279_ _280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_706_ _341_ _342_ _343_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_499_ _064_ net1 _155_ _156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_568_ _175_ _216_ _217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__527__A1 _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_353_ _042_ Datapath.i\[1\] _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_422_ Datapath.k\[2\] _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xinput8 co[1] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_405_ Datapath.k\[11\] _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 co[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__654__A3 _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_670_ Datapath.k\[16\] Datapath.k\[15\] _311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__590__A2 _237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__712__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__572__A2 _220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_653_ _290_ _291_ _294_ _295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_722_ _015_ clknet_2_2__leaf_clk Datapath.i\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_584_ Datapath.k\[9\] Datapath.k\[8\] _232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__735__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_705_ _047_ Datapath.k\[19\] _343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_567_ _214_ _215_ _216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_636_ _263_ _271_ _279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__536__A2 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_498_ _060_ Datapath.k\[0\] _037_ _155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__472__A1 _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__527__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_421_ Datapath.k\[3\] _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_41_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__518__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_352_ _041_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_14_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 co[2] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__454__A1 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_619_ _261_ _262_ _263_ _264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__509__A2 _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__445__A1 _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_404_ Datapath.k\[19\] Datapath.k\[18\] _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__675__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__427__A1 _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__469__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__657__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 co[5] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__646__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__639__A1 _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__501__I _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__392__B _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_652_ _293_ _294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_721_ _014_ clknet_2_3__leaf_clk Datapath.i\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_583_ _227_ _224_ _231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__539__B1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input10_I co[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__406__I Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_704_ _335_ _331_ _339_ _342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__481__A2 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_635_ _257_ _259_ _277_ _278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_566_ _198_ _207_ _215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_497_ _153_ _154_ _121_ _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input2_I co[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__472__A2 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__725__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_420_ _093_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_351_ _039_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__454__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_618_ Datapath.k\[12\] Datapath.k\[11\] _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_549_ _194_ _198_ _200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__445__A2 _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_403_ _075_ _076_ _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__372__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__427__A2 _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__675__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__363__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__666__A2 _279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__418__A2 _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__414__I Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__657__A2 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput13 co[6] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__584__A1 Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__639__A2 _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__575__A1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__409__I Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_720_ _013_ clknet_2_2__leaf_clk Datapath.i\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_651_ _090_ _292_ _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_582_ _229_ _230_ _076_ _158_ _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__539__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__539__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__422__I Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_634_ _265_ _272_ _277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_703_ _340_ _317_ _341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__481__A3 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__744__D FSM.NS\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_496_ _149_ _059_ _058_ _154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_565_ _188_ _179_ _214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__472__A3 _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__417__I _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_350_ net18 _040_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_617_ _099_ _079_ _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_479_ _134_ _138_ _141_ _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_548_ _194_ _198_ _199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__678__B1 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_402_ Datapath.k\[8\] _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__372__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__427__A3 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__363__A2 Datapath.i\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__715__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__418__A3 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput14 co[7] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_14_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__738__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__584__A2 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__425__I Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__575__A2 Datapath.k\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_650_ Datapath.k\[15\] Datapath.k\[14\] _292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_581_ net15 _120_ Datapath.k\[9\] _102_ _046_ _230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_16_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__484__A1 _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_633_ _275_ _276_ _098_ _047_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_702_ _335_ _331_ _339_ _340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_495_ _152_ Datapath.i\[15\] _153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_564_ _211_ _212_ _213_ _158_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__457__A1 _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__679__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__620__A1 _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__439__A1 _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_616_ _260_ _261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_547_ _196_ _197_ _198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_478_ _140_ _141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__678__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__678__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__602__A1 Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__428__I _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_401_ Datapath.k\[9\] _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__427__A4 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__520__B1 _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput15 co[8] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__502__B1 _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__531__I Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__687__B _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__616__I _260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__351__I _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__728__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__493__A2 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_580_ _227_ _064_ _228_ _229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__484__A2 Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__346__I _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__475__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_563_ Datapath.k\[7\] _213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_632_ Datapath.k\[14\] _103_ _038_ net5 _046_ _276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_701_ _078_ _338_ _339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_494_ _151_ _152_ _121_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_5_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__448__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__620__A2 _263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__384__A1 _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__589__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_615_ _257_ _259_ _260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_546_ Datapath.k\[6\] Datapath.k\[5\] _197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_477_ _139_ Datapath.i\[10\] _140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__678__A2 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__602__A2 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__534__I Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__366__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_400_ _072_ _039_ _073_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_529_ _180_ _064_ _181_ _182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__354__I _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__520__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 co[9] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__502__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__452__I _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__705__A1 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__632__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_700_ Datapath.k\[19\] Datapath.k\[18\] _338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__623__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_631_ _273_ _274_ _036_ _275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_562_ net14 _120_ Datapath.k\[8\] _102_ _046_ _212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_493_ _149_ _058_ _152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__357__I Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__718__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_614_ _258_ _242_ _248_ _259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_476_ _138_ _139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_545_ _195_ _196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__366__A2 _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__596__A2 _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_459_ _125_ Datapath.i\[6\] _062_ _126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_528_ _175_ _179_ _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__511__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__502__A2 _157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 st net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__650__A1 Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__632__A1 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__623__A1 Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_630_ _270_ _272_ _274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_492_ _149_ _058_ _151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_561_ _208_ _064_ _210_ _211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_613_ _255_ _239_ _258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_475_ _135_ _037_ _123_ _137_ _138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_544_ Datapath.k\[6\] Datapath.k\[5\] _195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__708__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_527_ _175_ _179_ _180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_389_ _036_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_458_ _119_ _121_ _125_ _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__505__B1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__511__A3 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__487__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__411__A2 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__650__A2 Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__469__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__641__A2 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__396__A1 _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__632__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__623__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_560_ _200_ _195_ _209_ _210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__741__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_491_ _150_ _121_ _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__378__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__614__A2 _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_689_ Datapath.k\[17\] Datapath.k\[15\] Datapath.k\[16\] _328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__605__A2 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_543_ _181_ _193_ _087_ _194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_612_ _217_ _220_ _256_ _257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_474_ _136_ _137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__474__I _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__532__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__649__I _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__523__A1 Datapath.k\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__514__A1 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_526_ _177_ _178_ _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__505__B2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_457_ _113_ _124_ _125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_388_ _047_ net17 _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__600__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_509_ _163_ _086_ _164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__505__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__521__B Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__496__A3 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input17_I st vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input9_I co[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__387__I _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__608__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_490_ Datapath.i\[13\] _146_ _149_ _150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__614__A3 _248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_688_ _314_ _084_ _321_ _327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__541__A2 _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_473_ Datapath.i\[9\] Datapath.i\[8\] _136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_542_ _192_ _193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_611_ _238_ _255_ _256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__599__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__523__A2 Datapath.k\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__731__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__514__A2 Datapath.k\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_525_ Datapath.k\[4\] Datapath.k\[3\] _178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_456_ _123_ _124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__505__A2 _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_387_ _061_ _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__441__A1 _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__432__A1 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__499__A1 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__423__A1 _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_508_ _161_ _162_ _163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_439_ _106_ _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__562__B1 Datapath.k\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__617__A1 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__608__A1 Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_687_ _325_ _326_ _121_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__550__A3 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_610_ _243_ _249_ _255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_472_ _111_ _051_ _050_ _135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_541_ _186_ _095_ _184_ _192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_739_ _032_ clknet_2_3__leaf_clk Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_386_ _038_ _060_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_524_ _176_ _177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_455_ _122_ _045_ _123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__441__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__519__C _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__432__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__499__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__423__A2 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_438_ Datapath.i\[2\] _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__721__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_369_ Datapath.i\[8\] _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_507_ Datapath.k\[2\] Datapath.k\[1\] _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__350__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__653__A2 _291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__744__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__399__A1 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__626__A2 _262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__562__B2 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__617__A2 _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__553__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__608__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__543__B _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__544__A1 Datapath.k\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_686_ _042_ Datapath.k\[17\] Datapath.k\[18\] _060_ _326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_540_ _190_ _191_ _186_ _158_ _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_471_ _062_ Datapath.i\[10\] _134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__517__A1 _165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_738_ _031_ clknet_2_2__leaf_clk Datapath.k\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_669_ _083_ _088_ _310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__508__A1 _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_523_ Datapath.k\[4\] Datapath.k\[3\] _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_385_ FSM.CS\[0\] _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_9_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_454_ Datapath.i\[5\] Datapath.i\[4\] _122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__B1 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_506_ _096_ _065_ _161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_437_ _043_ _107_ _108_ _040_ _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_368_ net18 _051_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__647__B1 _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__350__A2 _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__580__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__399__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__711__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__734__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input15_I co[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__544__A2 Datapath.k\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_685_ _322_ _317_ _324_ _325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I co[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__471__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__517__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_470_ _053_ _131_ _133_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_737_ _030_ clknet_2_2__leaf_clk Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_599_ _244_ _064_ _245_ _246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_668_ _304_ _308_ _309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__508__A2 _162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__444__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__435__A1 _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_522_ _165_ _170_ _174_ _175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_453_ _120_ _121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_384_ _039_ _059_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__426__A1 _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__459__B _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__665__A1 _283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__551__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__656__A1 Datapath.k\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_505_ net9 _121_ Datapath.k\[3\] _103_ _042_ _160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_436_ Datapath.i\[1\] _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_367_ Datapath.i\[7\] _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__647__B2 _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__629__A1 _270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_419_ Datapath.k\[7\] Datapath.k\[6\] _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__401__I Datapath.k\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__480__A2 _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_684_ _315_ _311_ _323_ _324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__471__A2 Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__517__A3 _170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_736_ _029_ clknet_2_0__leaf_clk Datapath.k\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__724__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_667_ _305_ _307_ _308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_598_ _240_ _243_ _245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__692__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__444__A2 Datapath.i\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__380__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__435__A2 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_521_ Datapath.k\[3\] Datapath.k\[1\] Datapath.k\[2\] _174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_383_ Datapath.i\[15\] _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_452_ _061_ _120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_17_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__426__A2 _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_719_ _012_ clknet_2_2__leaf_clk Datapath.i\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__353__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__656__A2 _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_435_ _106_ _037_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_504_ _060_ _065_ _096_ _073_ _159_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_366_ net18 _050_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__562__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__629__A2 _272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__565__A1 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_349_ Datapath.i\[0\] _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_418_ _085_ _086_ _087_ _091_ _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__538__A1 _185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__701__A1 _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_683_ _084_ _321_ _323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_735_ _028_ clknet_2_0__leaf_clk Datapath.k\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_666_ _300_ _279_ _306_ _307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_597_ _240_ _243_ _244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__601__B1 _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_520_ _172_ _173_ _095_ _158_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_382_ _039_ _058_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_451_ _118_ Datapath.i\[5\] _119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_718_ _011_ clknet_2_2__leaf_clk Datapath.i\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_649_ _283_ _291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__714__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_503_ _121_ net8 _159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_434_ Datapath.i\[1\] Datapath.i\[0\] _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_365_ Datapath.i\[6\] _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__737__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__415__I Datapath.k\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__565__A2 _179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_348_ _039_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_417_ _090_ _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__483__A1 _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__538__A2 _188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__529__A2 _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_682_ _320_ _084_ _321_ _322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__465__A1 _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I co[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__686__A1 _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__686__B2 _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_665_ _283_ _292_ _306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_734_ _027_ clknet_2_1__leaf_clk Datapath.k\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_596_ _241_ _242_ _243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I co[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__601__B2 _158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_450_ _116_ _118_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_381_ Datapath.i\[14\] _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__581__C _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_717_ _010_ clknet_2_2__leaf_clk Datapath.i\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_648_ _278_ _280_ _284_ _290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_579_ _222_ _225_ _228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_433_ _039_ _040_ _105_ _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_502_ _156_ _157_ _086_ _158_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_364_ _049_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__587__B _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_416_ _088_ _089_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_347_ _036_ _038_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__492__A2 _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__727__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__529__A3 _181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_681_ Datapath.k\[17\] Datapath.k\[16\] _321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__392__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__447__A2 Datapath.i\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__686__A2 Datapath.k\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_664_ _259_ _302_ _305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_733_ _026_ clknet_2_1__leaf_clk Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_595_ Datapath.k\[10\] Datapath.k\[9\] _242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__524__I _176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_380_ net18 _057_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__659__A2 _293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 x[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_716_ _009_ clknet_2_2__leaf_clk Datapath.i\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__595__A1 Datapath.k\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_578_ _226_ _227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_647_ _288_ _289_ _089_ _047_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__347__A1 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

