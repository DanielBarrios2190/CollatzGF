magic
tech gf180mcuC
magscale 1 10
timestamp 1670117119
<< metal1 >>
rect 1344 40794 42560 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 42560 40794
rect 1344 40708 42560 40742
rect 1344 40010 42560 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 42560 40010
rect 1344 39924 42560 39958
rect 1344 39226 42560 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 42560 39226
rect 1344 39140 42560 39174
rect 1344 38442 42560 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 42560 38442
rect 1344 38356 42560 38390
rect 1344 37658 42560 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 42560 37658
rect 1344 37572 42560 37606
rect 1344 36874 42560 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 42560 36874
rect 1344 36788 42560 36822
rect 1344 36090 42560 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 42560 36090
rect 1344 36004 42560 36038
rect 1344 35306 42560 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 42560 35306
rect 1344 35220 42560 35254
rect 1344 34522 42560 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 42560 34522
rect 1344 34436 42560 34470
rect 1344 33738 42560 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 42560 33738
rect 1344 33652 42560 33686
rect 1344 32954 42560 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 42560 32954
rect 1344 32868 42560 32902
rect 1344 32170 42560 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 42560 32170
rect 1344 32084 42560 32118
rect 1344 31386 42560 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 42560 31386
rect 1344 31300 42560 31334
rect 1344 30602 42560 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 42560 30602
rect 1344 30516 42560 30550
rect 1344 29818 42560 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 42560 29818
rect 1344 29732 42560 29766
rect 1344 29034 42560 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 42560 29034
rect 1344 28948 42560 28982
rect 1344 28250 42560 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 42560 28250
rect 1344 28164 42560 28198
rect 1344 27466 42560 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 42560 27466
rect 1344 27380 42560 27414
rect 1344 26682 42560 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 42560 26682
rect 1344 26596 42560 26630
rect 1344 25898 42560 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 42560 25898
rect 1344 25812 42560 25846
rect 1344 25114 42560 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 42560 25114
rect 1344 25028 42560 25062
rect 30158 24610 30210 24622
rect 30158 24546 30210 24558
rect 30606 24610 30658 24622
rect 30606 24546 30658 24558
rect 31838 24610 31890 24622
rect 31838 24546 31890 24558
rect 41582 24610 41634 24622
rect 41582 24546 41634 24558
rect 1344 24330 42560 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 42560 24330
rect 1344 24244 42560 24278
rect 32050 24110 32062 24162
rect 32114 24159 32126 24162
rect 32946 24159 32958 24162
rect 32114 24113 32958 24159
rect 32114 24110 32126 24113
rect 32946 24110 32958 24113
rect 33010 24110 33022 24162
rect 28030 24050 28082 24062
rect 28030 23986 28082 23998
rect 30494 24050 30546 24062
rect 30494 23986 30546 23998
rect 32958 24050 33010 24062
rect 32958 23986 33010 23998
rect 35758 24050 35810 24062
rect 35758 23986 35810 23998
rect 36878 24050 36930 24062
rect 36878 23986 36930 23998
rect 34190 23938 34242 23950
rect 34190 23874 34242 23886
rect 39454 23826 39506 23838
rect 39454 23762 39506 23774
rect 28702 23714 28754 23726
rect 28702 23650 28754 23662
rect 29598 23714 29650 23726
rect 29598 23650 29650 23662
rect 30046 23714 30098 23726
rect 30046 23650 30098 23662
rect 31166 23714 31218 23726
rect 31166 23650 31218 23662
rect 31502 23714 31554 23726
rect 31502 23650 31554 23662
rect 32062 23714 32114 23726
rect 32062 23650 32114 23662
rect 32510 23714 32562 23726
rect 32510 23650 32562 23662
rect 33294 23714 33346 23726
rect 33294 23650 33346 23662
rect 33854 23714 33906 23726
rect 33854 23650 33906 23662
rect 35310 23714 35362 23726
rect 35310 23650 35362 23662
rect 36430 23714 36482 23726
rect 36430 23650 36482 23662
rect 37774 23714 37826 23726
rect 37774 23650 37826 23662
rect 38222 23714 38274 23726
rect 38222 23650 38274 23662
rect 38670 23714 38722 23726
rect 38670 23650 38722 23662
rect 39118 23714 39170 23726
rect 39118 23650 39170 23662
rect 40238 23714 40290 23726
rect 40238 23650 40290 23662
rect 40686 23714 40738 23726
rect 40686 23650 40738 23662
rect 41358 23714 41410 23726
rect 41358 23650 41410 23662
rect 41806 23714 41858 23726
rect 41806 23650 41858 23662
rect 1344 23546 42560 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 42560 23546
rect 1344 23460 42560 23494
rect 32958 23378 33010 23390
rect 32958 23314 33010 23326
rect 32510 23266 32562 23278
rect 32510 23202 32562 23214
rect 39678 23266 39730 23278
rect 39678 23202 39730 23214
rect 42030 23266 42082 23278
rect 42030 23202 42082 23214
rect 29710 23154 29762 23166
rect 29710 23090 29762 23102
rect 37662 23154 37714 23166
rect 37662 23090 37714 23102
rect 26238 23042 26290 23054
rect 26238 22978 26290 22990
rect 26574 23042 26626 23054
rect 26574 22978 26626 22990
rect 27134 23042 27186 23054
rect 27134 22978 27186 22990
rect 27582 23042 27634 23054
rect 27582 22978 27634 22990
rect 28254 23042 28306 23054
rect 28254 22978 28306 22990
rect 28590 23042 28642 23054
rect 28590 22978 28642 22990
rect 29374 23042 29426 23054
rect 29374 22978 29426 22990
rect 30494 23042 30546 23054
rect 30494 22978 30546 22990
rect 30830 23042 30882 23054
rect 30830 22978 30882 22990
rect 31614 23042 31666 23054
rect 31614 22978 31666 22990
rect 31950 23042 32002 23054
rect 31950 22978 32002 22990
rect 33518 23042 33570 23054
rect 33518 22978 33570 22990
rect 33966 23042 34018 23054
rect 33966 22978 34018 22990
rect 34526 23042 34578 23054
rect 34526 22978 34578 22990
rect 34862 23042 34914 23054
rect 34862 22978 34914 22990
rect 35422 23042 35474 23054
rect 35422 22978 35474 22990
rect 35870 23042 35922 23054
rect 35870 22978 35922 22990
rect 36206 23042 36258 23054
rect 36206 22978 36258 22990
rect 36766 23042 36818 23054
rect 36766 22978 36818 22990
rect 37102 23042 37154 23054
rect 37102 22978 37154 22990
rect 38334 23042 38386 23054
rect 38334 22978 38386 22990
rect 38782 23042 38834 23054
rect 38782 22978 38834 22990
rect 39230 23042 39282 23054
rect 39230 22978 39282 22990
rect 40238 23042 40290 23054
rect 40238 22978 40290 22990
rect 40686 23042 40738 23054
rect 40686 22978 40738 22990
rect 41470 23042 41522 23054
rect 41470 22978 41522 22990
rect 35634 22878 35646 22930
rect 35698 22927 35710 22930
rect 36754 22927 36766 22930
rect 35698 22881 36766 22927
rect 35698 22878 35710 22881
rect 36754 22878 36766 22881
rect 36818 22878 36830 22930
rect 1344 22762 42560 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 42560 22762
rect 1344 22676 42560 22710
rect 35970 22542 35982 22594
rect 36034 22591 36046 22594
rect 36418 22591 36430 22594
rect 36034 22545 36430 22591
rect 36034 22542 36046 22545
rect 36418 22542 36430 22545
rect 36482 22542 36494 22594
rect 24782 22482 24834 22494
rect 3266 22430 3278 22482
rect 3330 22430 3342 22482
rect 24782 22418 24834 22430
rect 25230 22482 25282 22494
rect 25230 22418 25282 22430
rect 25566 22482 25618 22494
rect 25566 22418 25618 22430
rect 26014 22482 26066 22494
rect 26014 22418 26066 22430
rect 26462 22482 26514 22494
rect 26462 22418 26514 22430
rect 29486 22482 29538 22494
rect 29486 22418 29538 22430
rect 30046 22482 30098 22494
rect 30046 22418 30098 22430
rect 31390 22482 31442 22494
rect 31390 22418 31442 22430
rect 31726 22482 31778 22494
rect 31726 22418 31778 22430
rect 32174 22482 32226 22494
rect 32174 22418 32226 22430
rect 32622 22482 32674 22494
rect 32622 22418 32674 22430
rect 34190 22482 34242 22494
rect 34190 22418 34242 22430
rect 35086 22482 35138 22494
rect 35086 22418 35138 22430
rect 36430 22482 36482 22494
rect 38546 22430 38558 22482
rect 38610 22479 38622 22482
rect 38882 22479 38894 22482
rect 38610 22433 38894 22479
rect 38610 22430 38622 22433
rect 38882 22430 38894 22433
rect 38946 22430 38958 22482
rect 36430 22418 36482 22430
rect 30494 22370 30546 22382
rect 30494 22306 30546 22318
rect 37886 22370 37938 22382
rect 38882 22318 38894 22370
rect 38946 22318 38958 22370
rect 37886 22306 37938 22318
rect 27806 22258 27858 22270
rect 1922 22206 1934 22258
rect 1986 22206 1998 22258
rect 27806 22194 27858 22206
rect 38334 22258 38386 22270
rect 40002 22206 40014 22258
rect 40066 22206 40078 22258
rect 38334 22194 38386 22206
rect 26910 22146 26962 22158
rect 26910 22082 26962 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 30942 22146 30994 22158
rect 30942 22082 30994 22094
rect 33406 22146 33458 22158
rect 33406 22082 33458 22094
rect 33742 22146 33794 22158
rect 33742 22082 33794 22094
rect 34750 22146 34802 22158
rect 34750 22082 34802 22094
rect 35534 22146 35586 22158
rect 35534 22082 35586 22094
rect 35982 22146 36034 22158
rect 35982 22082 36034 22094
rect 37438 22146 37490 22158
rect 37438 22082 37490 22094
rect 40574 22146 40626 22158
rect 40574 22082 40626 22094
rect 41022 22146 41074 22158
rect 41022 22082 41074 22094
rect 41694 22146 41746 22158
rect 41694 22082 41746 22094
rect 42030 22146 42082 22158
rect 42030 22082 42082 22094
rect 1344 21978 42560 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 42560 21978
rect 1344 21892 42560 21926
rect 1822 21810 1874 21822
rect 1822 21746 1874 21758
rect 28814 21810 28866 21822
rect 28814 21746 28866 21758
rect 32174 21810 32226 21822
rect 32174 21746 32226 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 35758 21810 35810 21822
rect 35758 21746 35810 21758
rect 37550 21810 37602 21822
rect 37550 21746 37602 21758
rect 38894 21810 38946 21822
rect 38894 21746 38946 21758
rect 42030 21810 42082 21822
rect 42030 21746 42082 21758
rect 26686 21586 26738 21598
rect 26686 21522 26738 21534
rect 34078 21586 34130 21598
rect 34078 21522 34130 21534
rect 24110 21474 24162 21486
rect 24110 21410 24162 21422
rect 24558 21474 24610 21486
rect 24558 21410 24610 21422
rect 24894 21474 24946 21486
rect 24894 21410 24946 21422
rect 25566 21474 25618 21486
rect 25566 21410 25618 21422
rect 26238 21474 26290 21486
rect 26238 21410 26290 21422
rect 27134 21474 27186 21486
rect 27134 21410 27186 21422
rect 27582 21474 27634 21486
rect 27582 21410 27634 21422
rect 28030 21474 28082 21486
rect 28030 21410 28082 21422
rect 28478 21474 28530 21486
rect 28478 21410 28530 21422
rect 29262 21474 29314 21486
rect 29262 21410 29314 21422
rect 30158 21474 30210 21486
rect 30158 21410 30210 21422
rect 30494 21474 30546 21486
rect 30494 21410 30546 21422
rect 31054 21474 31106 21486
rect 31054 21410 31106 21422
rect 31726 21474 31778 21486
rect 31726 21410 31778 21422
rect 32734 21474 32786 21486
rect 32734 21410 32786 21422
rect 33630 21474 33682 21486
rect 33630 21410 33682 21422
rect 34414 21474 34466 21486
rect 34414 21410 34466 21422
rect 35422 21474 35474 21486
rect 35422 21410 35474 21422
rect 36318 21474 36370 21486
rect 36318 21410 36370 21422
rect 36766 21474 36818 21486
rect 36766 21410 36818 21422
rect 37214 21474 37266 21486
rect 37214 21410 37266 21422
rect 37998 21474 38050 21486
rect 37998 21410 38050 21422
rect 38446 21474 38498 21486
rect 38446 21410 38498 21422
rect 39342 21474 39394 21486
rect 39342 21410 39394 21422
rect 40014 21474 40066 21486
rect 40014 21410 40066 21422
rect 40462 21474 40514 21486
rect 40462 21410 40514 21422
rect 41470 21474 41522 21486
rect 41470 21410 41522 21422
rect 37202 21310 37214 21362
rect 37266 21359 37278 21362
rect 38098 21359 38110 21362
rect 37266 21313 38110 21359
rect 37266 21310 37278 21313
rect 38098 21310 38110 21313
rect 38162 21310 38174 21362
rect 1344 21194 42560 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 42560 21194
rect 1344 21108 42560 21142
rect 33506 20974 33518 21026
rect 33570 21023 33582 21026
rect 34402 21023 34414 21026
rect 33570 20977 34414 21023
rect 33570 20974 33582 20977
rect 34402 20974 34414 20977
rect 34466 21023 34478 21026
rect 34850 21023 34862 21026
rect 34466 20977 34862 21023
rect 34466 20974 34478 20977
rect 34850 20974 34862 20977
rect 34914 21023 34926 21026
rect 35074 21023 35086 21026
rect 34914 20977 35086 21023
rect 34914 20974 34926 20977
rect 35074 20974 35086 20977
rect 35138 20974 35150 21026
rect 35298 20974 35310 21026
rect 35362 21023 35374 21026
rect 36194 21023 36206 21026
rect 35362 20977 36206 21023
rect 35362 20974 35374 20977
rect 36194 20974 36206 20977
rect 36258 20974 36270 21026
rect 22990 20914 23042 20926
rect 22990 20850 23042 20862
rect 23438 20914 23490 20926
rect 23438 20850 23490 20862
rect 23886 20914 23938 20926
rect 23886 20850 23938 20862
rect 29934 20914 29986 20926
rect 29934 20850 29986 20862
rect 31278 20914 31330 20926
rect 31278 20850 31330 20862
rect 32622 20914 32674 20926
rect 32622 20850 32674 20862
rect 33070 20914 33122 20926
rect 33070 20850 33122 20862
rect 33518 20914 33570 20926
rect 33518 20850 33570 20862
rect 34414 20914 34466 20926
rect 34414 20850 34466 20862
rect 34862 20914 34914 20926
rect 34862 20850 34914 20862
rect 35310 20914 35362 20926
rect 35310 20850 35362 20862
rect 35758 20914 35810 20926
rect 35758 20850 35810 20862
rect 38782 20914 38834 20926
rect 38782 20850 38834 20862
rect 41246 20914 41298 20926
rect 41246 20850 41298 20862
rect 42030 20914 42082 20926
rect 42030 20850 42082 20862
rect 26238 20802 26290 20814
rect 26238 20738 26290 20750
rect 36206 20802 36258 20814
rect 36206 20738 36258 20750
rect 37438 20802 37490 20814
rect 37438 20738 37490 20750
rect 24334 20690 24386 20702
rect 24334 20626 24386 20638
rect 26574 20690 26626 20702
rect 26574 20626 26626 20638
rect 28702 20690 28754 20702
rect 28702 20626 28754 20638
rect 36654 20690 36706 20702
rect 36654 20626 36706 20638
rect 24670 20578 24722 20590
rect 24670 20514 24722 20526
rect 25230 20578 25282 20590
rect 25230 20514 25282 20526
rect 25790 20578 25842 20590
rect 25790 20514 25842 20526
rect 27022 20578 27074 20590
rect 27022 20514 27074 20526
rect 27918 20578 27970 20590
rect 27918 20514 27970 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 29486 20578 29538 20590
rect 29486 20514 29538 20526
rect 30494 20578 30546 20590
rect 30494 20514 30546 20526
rect 30942 20578 30994 20590
rect 30942 20514 30994 20526
rect 31838 20578 31890 20590
rect 31838 20514 31890 20526
rect 32286 20578 32338 20590
rect 32286 20514 32338 20526
rect 33966 20578 34018 20590
rect 33966 20514 34018 20526
rect 37886 20578 37938 20590
rect 37886 20514 37938 20526
rect 38334 20578 38386 20590
rect 38334 20514 38386 20526
rect 39230 20578 39282 20590
rect 39230 20514 39282 20526
rect 40014 20578 40066 20590
rect 40014 20514 40066 20526
rect 40462 20578 40514 20590
rect 40462 20514 40514 20526
rect 1344 20410 42560 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 42560 20410
rect 1344 20324 42560 20358
rect 31838 20242 31890 20254
rect 31838 20178 31890 20190
rect 34862 20242 34914 20254
rect 34862 20178 34914 20190
rect 22878 20130 22930 20142
rect 22878 20066 22930 20078
rect 23326 20130 23378 20142
rect 23326 20066 23378 20078
rect 25566 20130 25618 20142
rect 25566 20066 25618 20078
rect 39342 20130 39394 20142
rect 39342 20066 39394 20078
rect 26014 20018 26066 20030
rect 26014 19954 26066 19966
rect 27806 20018 27858 20030
rect 27806 19954 27858 19966
rect 33518 20018 33570 20030
rect 33518 19954 33570 19966
rect 34414 20018 34466 20030
rect 34414 19954 34466 19966
rect 37998 20018 38050 20030
rect 37998 19954 38050 19966
rect 22094 19906 22146 19918
rect 22094 19842 22146 19854
rect 22542 19906 22594 19918
rect 22542 19842 22594 19854
rect 23886 19906 23938 19918
rect 23886 19842 23938 19854
rect 24222 19906 24274 19918
rect 24222 19842 24274 19854
rect 24670 19906 24722 19918
rect 24670 19842 24722 19854
rect 26574 19906 26626 19918
rect 26574 19842 26626 19854
rect 26910 19906 26962 19918
rect 26910 19842 26962 19854
rect 27470 19906 27522 19918
rect 27470 19842 27522 19854
rect 28254 19906 28306 19918
rect 28254 19842 28306 19854
rect 28702 19906 28754 19918
rect 28702 19842 28754 19854
rect 29262 19906 29314 19918
rect 29262 19842 29314 19854
rect 29598 19906 29650 19918
rect 29598 19842 29650 19854
rect 30158 19906 30210 19918
rect 30158 19842 30210 19854
rect 30494 19906 30546 19918
rect 30494 19842 30546 19854
rect 31054 19906 31106 19918
rect 31054 19842 31106 19854
rect 31390 19906 31442 19918
rect 31390 19842 31442 19854
rect 32286 19906 32338 19918
rect 32286 19842 32338 19854
rect 32846 19906 32898 19918
rect 32846 19842 32898 19854
rect 33966 19906 34018 19918
rect 33966 19842 34018 19854
rect 35422 19906 35474 19918
rect 35422 19842 35474 19854
rect 35758 19906 35810 19918
rect 35758 19842 35810 19854
rect 36206 19906 36258 19918
rect 36206 19842 36258 19854
rect 36766 19906 36818 19918
rect 36766 19842 36818 19854
rect 37102 19906 37154 19918
rect 37102 19842 37154 19854
rect 37550 19906 37602 19918
rect 37550 19842 37602 19854
rect 38446 19906 38498 19918
rect 38446 19842 38498 19854
rect 38894 19906 38946 19918
rect 38894 19842 38946 19854
rect 39790 19906 39842 19918
rect 39790 19842 39842 19854
rect 40350 19906 40402 19918
rect 40350 19842 40402 19854
rect 40798 19906 40850 19918
rect 40798 19842 40850 19854
rect 41470 19906 41522 19918
rect 41470 19842 41522 19854
rect 41918 19906 41970 19918
rect 41918 19842 41970 19854
rect 21970 19742 21982 19794
rect 22034 19791 22046 19794
rect 23314 19791 23326 19794
rect 22034 19745 23326 19791
rect 22034 19742 22046 19745
rect 23314 19742 23326 19745
rect 23378 19742 23390 19794
rect 28690 19742 28702 19794
rect 28754 19791 28766 19794
rect 29474 19791 29486 19794
rect 28754 19745 29486 19791
rect 28754 19742 28766 19745
rect 29474 19742 29486 19745
rect 29538 19742 29550 19794
rect 37314 19742 37326 19794
rect 37378 19791 37390 19794
rect 37874 19791 37886 19794
rect 37378 19745 37886 19791
rect 37378 19742 37390 19745
rect 37874 19742 37886 19745
rect 37938 19742 37950 19794
rect 1344 19626 42560 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 42560 19626
rect 1344 19540 42560 19574
rect 37426 19406 37438 19458
rect 37490 19455 37502 19458
rect 38322 19455 38334 19458
rect 37490 19409 38334 19455
rect 37490 19406 37502 19409
rect 38322 19406 38334 19409
rect 38386 19406 38398 19458
rect 39666 19406 39678 19458
rect 39730 19455 39742 19458
rect 40226 19455 40238 19458
rect 39730 19409 40238 19455
rect 39730 19406 39742 19409
rect 40226 19406 40238 19409
rect 40290 19406 40302 19458
rect 41234 19406 41246 19458
rect 41298 19455 41310 19458
rect 41906 19455 41918 19458
rect 41298 19409 41918 19455
rect 41298 19406 41310 19409
rect 41906 19406 41918 19409
rect 41970 19406 41982 19458
rect 21646 19346 21698 19358
rect 21646 19282 21698 19294
rect 27694 19346 27746 19358
rect 27694 19282 27746 19294
rect 28590 19346 28642 19358
rect 28590 19282 28642 19294
rect 33630 19346 33682 19358
rect 33630 19282 33682 19294
rect 35086 19346 35138 19358
rect 35086 19282 35138 19294
rect 37886 19346 37938 19358
rect 37886 19282 37938 19294
rect 40238 19346 40290 19358
rect 40238 19282 40290 19294
rect 42030 19346 42082 19358
rect 42030 19282 42082 19294
rect 23326 19234 23378 19246
rect 23326 19170 23378 19182
rect 23662 19234 23714 19246
rect 34190 19234 34242 19246
rect 25218 19182 25230 19234
rect 25282 19182 25294 19234
rect 23662 19170 23714 19182
rect 34190 19170 34242 19182
rect 25006 19122 25058 19134
rect 25006 19058 25058 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 26238 19122 26290 19134
rect 26238 19058 26290 19070
rect 39678 19122 39730 19134
rect 39678 19058 39730 19070
rect 20862 19010 20914 19022
rect 20862 18946 20914 18958
rect 22094 19010 22146 19022
rect 22094 18946 22146 18958
rect 22542 19010 22594 19022
rect 22542 18946 22594 18958
rect 22990 19010 23042 19022
rect 22990 18946 23042 18958
rect 23550 19010 23602 19022
rect 23550 18946 23602 18958
rect 24110 19010 24162 19022
rect 24110 18946 24162 18958
rect 25454 19010 25506 19022
rect 25454 18946 25506 18958
rect 25566 19010 25618 19022
rect 25566 18946 25618 18958
rect 26126 19010 26178 19022
rect 26126 18946 26178 18958
rect 26686 19010 26738 19022
rect 26686 18946 26738 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 28142 19010 28194 19022
rect 28142 18946 28194 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 29934 19010 29986 19022
rect 29934 18946 29986 18958
rect 30718 19010 30770 19022
rect 30718 18946 30770 18958
rect 31166 19010 31218 19022
rect 31166 18946 31218 18958
rect 31614 19010 31666 19022
rect 31614 18946 31666 18958
rect 32286 19010 32338 19022
rect 32286 18946 32338 18958
rect 32846 19010 32898 19022
rect 32846 18946 32898 18958
rect 33294 19010 33346 19022
rect 33294 18946 33346 18958
rect 34638 19010 34690 19022
rect 34638 18946 34690 18958
rect 35758 19010 35810 19022
rect 35758 18946 35810 18958
rect 36206 19010 36258 19022
rect 36206 18946 36258 18958
rect 36654 19010 36706 19022
rect 36654 18946 36706 18958
rect 37438 19010 37490 19022
rect 37438 18946 37490 18958
rect 38334 19010 38386 19022
rect 38334 18946 38386 18958
rect 38782 19010 38834 19022
rect 38782 18946 38834 18958
rect 39230 19010 39282 19022
rect 39230 18946 39282 18958
rect 40686 19010 40738 19022
rect 40686 18946 40738 18958
rect 41246 19010 41298 19022
rect 41246 18946 41298 18958
rect 41694 19010 41746 19022
rect 41694 18946 41746 18958
rect 1344 18842 42560 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 42560 18842
rect 1344 18756 42560 18790
rect 24110 18674 24162 18686
rect 24110 18610 24162 18622
rect 29822 18674 29874 18686
rect 29822 18610 29874 18622
rect 24334 18562 24386 18574
rect 24334 18498 24386 18510
rect 23886 18450 23938 18462
rect 20626 18398 20638 18450
rect 20690 18398 20702 18450
rect 23886 18386 23938 18398
rect 24446 18450 24498 18462
rect 29934 18450 29986 18462
rect 39006 18450 39058 18462
rect 26114 18398 26126 18450
rect 26178 18398 26190 18450
rect 36082 18398 36094 18450
rect 36146 18447 36158 18450
rect 36306 18447 36318 18450
rect 36146 18401 36318 18447
rect 36146 18398 36158 18401
rect 36306 18398 36318 18401
rect 36370 18398 36382 18450
rect 24446 18386 24498 18398
rect 29934 18386 29986 18398
rect 39006 18386 39058 18398
rect 39454 18450 39506 18462
rect 39454 18386 39506 18398
rect 41918 18450 41970 18462
rect 41918 18386 41970 18398
rect 20078 18338 20130 18350
rect 30606 18338 30658 18350
rect 21298 18286 21310 18338
rect 21362 18286 21374 18338
rect 23426 18286 23438 18338
rect 23490 18286 23502 18338
rect 26786 18286 26798 18338
rect 26850 18286 26862 18338
rect 28914 18286 28926 18338
rect 28978 18286 28990 18338
rect 20078 18274 20130 18286
rect 30606 18274 30658 18286
rect 31054 18338 31106 18350
rect 31054 18274 31106 18286
rect 31502 18338 31554 18350
rect 31502 18274 31554 18286
rect 31950 18338 32002 18350
rect 31950 18274 32002 18286
rect 32398 18338 32450 18350
rect 32398 18274 32450 18286
rect 32958 18338 33010 18350
rect 32958 18274 33010 18286
rect 33518 18338 33570 18350
rect 33518 18274 33570 18286
rect 34078 18338 34130 18350
rect 34078 18274 34130 18286
rect 34862 18338 34914 18350
rect 34862 18274 34914 18286
rect 35422 18338 35474 18350
rect 35422 18274 35474 18286
rect 35870 18338 35922 18350
rect 35870 18274 35922 18286
rect 36430 18338 36482 18350
rect 36430 18274 36482 18286
rect 37102 18338 37154 18350
rect 37102 18274 37154 18286
rect 37662 18338 37714 18350
rect 37662 18274 37714 18286
rect 38110 18338 38162 18350
rect 38110 18274 38162 18286
rect 38558 18338 38610 18350
rect 38558 18274 38610 18286
rect 39902 18338 39954 18350
rect 39902 18274 39954 18286
rect 40462 18338 40514 18350
rect 40462 18274 40514 18286
rect 40798 18338 40850 18350
rect 40798 18274 40850 18286
rect 42030 18338 42082 18350
rect 42030 18274 42082 18286
rect 29822 18226 29874 18238
rect 29822 18162 29874 18174
rect 30494 18226 30546 18238
rect 30494 18162 30546 18174
rect 34974 18226 35026 18238
rect 36542 18226 36594 18238
rect 35522 18174 35534 18226
rect 35586 18223 35598 18226
rect 35858 18223 35870 18226
rect 35586 18177 35870 18223
rect 35586 18174 35598 18177
rect 35858 18174 35870 18177
rect 35922 18174 35934 18226
rect 34974 18162 35026 18174
rect 36542 18162 36594 18174
rect 37214 18226 37266 18238
rect 37874 18174 37886 18226
rect 37938 18223 37950 18226
rect 38546 18223 38558 18226
rect 37938 18177 38558 18223
rect 37938 18174 37950 18177
rect 38546 18174 38558 18177
rect 38610 18174 38622 18226
rect 40338 18174 40350 18226
rect 40402 18223 40414 18226
rect 40786 18223 40798 18226
rect 40402 18177 40798 18223
rect 40402 18174 40414 18177
rect 40786 18174 40798 18177
rect 40850 18174 40862 18226
rect 37214 18162 37266 18174
rect 1344 18058 42560 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 42560 18058
rect 1344 17972 42560 18006
rect 23438 17890 23490 17902
rect 23438 17826 23490 17838
rect 24782 17890 24834 17902
rect 24782 17826 24834 17838
rect 25454 17890 25506 17902
rect 25454 17826 25506 17838
rect 25790 17890 25842 17902
rect 25790 17826 25842 17838
rect 27358 17890 27410 17902
rect 27358 17826 27410 17838
rect 28142 17890 28194 17902
rect 28142 17826 28194 17838
rect 41246 17890 41298 17902
rect 41246 17826 41298 17838
rect 42030 17890 42082 17902
rect 42030 17826 42082 17838
rect 18622 17778 18674 17790
rect 18622 17714 18674 17726
rect 19070 17778 19122 17790
rect 19070 17714 19122 17726
rect 19854 17778 19906 17790
rect 19854 17714 19906 17726
rect 20862 17778 20914 17790
rect 20862 17714 20914 17726
rect 21758 17778 21810 17790
rect 21758 17714 21810 17726
rect 26014 17778 26066 17790
rect 26014 17714 26066 17726
rect 28590 17778 28642 17790
rect 28590 17714 28642 17726
rect 30942 17778 30994 17790
rect 41358 17778 41410 17790
rect 35298 17726 35310 17778
rect 35362 17726 35374 17778
rect 30942 17714 30994 17726
rect 41358 17714 41410 17726
rect 41918 17778 41970 17790
rect 41918 17714 41970 17726
rect 21646 17666 21698 17678
rect 21646 17602 21698 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 22318 17666 22370 17678
rect 24110 17666 24162 17678
rect 23762 17614 23774 17666
rect 23826 17614 23838 17666
rect 22318 17602 22370 17614
rect 24110 17602 24162 17614
rect 30046 17666 30098 17678
rect 30046 17602 30098 17614
rect 30270 17666 30322 17678
rect 38782 17666 38834 17678
rect 32498 17614 32510 17666
rect 32562 17614 32574 17666
rect 30270 17602 30322 17614
rect 38782 17602 38834 17614
rect 23550 17554 23602 17566
rect 23550 17490 23602 17502
rect 24894 17554 24946 17566
rect 24894 17490 24946 17502
rect 26574 17554 26626 17566
rect 26574 17490 26626 17502
rect 26910 17554 26962 17566
rect 26910 17490 26962 17502
rect 27470 17554 27522 17566
rect 27470 17490 27522 17502
rect 28030 17554 28082 17566
rect 28030 17490 28082 17502
rect 31054 17554 31106 17566
rect 35982 17554 36034 17566
rect 33170 17502 33182 17554
rect 33234 17502 33246 17554
rect 31054 17490 31106 17502
rect 35982 17490 36034 17502
rect 37550 17554 37602 17566
rect 37550 17490 37602 17502
rect 39230 17554 39282 17566
rect 39230 17490 39282 17502
rect 40574 17554 40626 17566
rect 40574 17490 40626 17502
rect 19518 17442 19570 17454
rect 19518 17378 19570 17390
rect 20414 17442 20466 17454
rect 20414 17378 20466 17390
rect 22990 17442 23042 17454
rect 22990 17378 23042 17390
rect 24782 17442 24834 17454
rect 24782 17378 24834 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 29822 17442 29874 17454
rect 29822 17378 29874 17390
rect 30158 17442 30210 17454
rect 30158 17378 30210 17390
rect 30830 17442 30882 17454
rect 30830 17378 30882 17390
rect 31278 17442 31330 17454
rect 31278 17378 31330 17390
rect 31838 17442 31890 17454
rect 31838 17378 31890 17390
rect 36094 17442 36146 17454
rect 36094 17378 36146 17390
rect 36318 17442 36370 17454
rect 36318 17378 36370 17390
rect 36654 17442 36706 17454
rect 36654 17378 36706 17390
rect 37662 17442 37714 17454
rect 37662 17378 37714 17390
rect 38110 17442 38162 17454
rect 38110 17378 38162 17390
rect 38222 17442 38274 17454
rect 38222 17378 38274 17390
rect 38446 17442 38498 17454
rect 38446 17378 38498 17390
rect 39342 17442 39394 17454
rect 39342 17378 39394 17390
rect 40014 17442 40066 17454
rect 40014 17378 40066 17390
rect 40686 17442 40738 17454
rect 40686 17378 40738 17390
rect 1344 17274 42560 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 42560 17274
rect 1344 17188 42560 17222
rect 18734 17106 18786 17118
rect 18734 17042 18786 17054
rect 19518 17106 19570 17118
rect 19518 17042 19570 17054
rect 19966 17106 20018 17118
rect 19966 17042 20018 17054
rect 21310 17106 21362 17118
rect 21310 17042 21362 17054
rect 23102 17106 23154 17118
rect 23102 17042 23154 17054
rect 24446 17106 24498 17118
rect 31614 17106 31666 17118
rect 26226 17054 26238 17106
rect 26290 17054 26302 17106
rect 24446 17042 24498 17054
rect 31614 17042 31666 17054
rect 32174 17106 32226 17118
rect 32174 17042 32226 17054
rect 37102 17106 37154 17118
rect 37102 17042 37154 17054
rect 37326 17106 37378 17118
rect 37326 17042 37378 17054
rect 38670 17106 38722 17118
rect 38670 17042 38722 17054
rect 21758 16994 21810 17006
rect 21758 16930 21810 16942
rect 23326 16994 23378 17006
rect 23326 16930 23378 16942
rect 23438 16994 23490 17006
rect 23438 16930 23490 16942
rect 24222 16994 24274 17006
rect 24222 16930 24274 16942
rect 30942 16994 30994 17006
rect 30942 16930 30994 16942
rect 31390 16994 31442 17006
rect 31390 16930 31442 16942
rect 31726 16994 31778 17006
rect 31726 16930 31778 16942
rect 32398 16994 32450 17006
rect 32398 16930 32450 16942
rect 38334 16994 38386 17006
rect 38334 16930 38386 16942
rect 39566 16994 39618 17006
rect 39566 16930 39618 16942
rect 40574 16994 40626 17006
rect 40574 16930 40626 16942
rect 41806 16994 41858 17006
rect 41806 16930 41858 16942
rect 41918 16994 41970 17006
rect 41918 16930 41970 16942
rect 15262 16882 15314 16894
rect 15262 16818 15314 16830
rect 17614 16882 17666 16894
rect 17614 16818 17666 16830
rect 18286 16882 18338 16894
rect 18286 16818 18338 16830
rect 20414 16882 20466 16894
rect 20414 16818 20466 16830
rect 20862 16882 20914 16894
rect 20862 16818 20914 16830
rect 22206 16882 22258 16894
rect 22206 16818 22258 16830
rect 22654 16882 22706 16894
rect 22654 16818 22706 16830
rect 24110 16882 24162 16894
rect 24110 16818 24162 16830
rect 24894 16882 24946 16894
rect 30382 16882 30434 16894
rect 32510 16882 32562 16894
rect 38558 16882 38610 16894
rect 27010 16830 27022 16882
rect 27074 16830 27086 16882
rect 30706 16830 30718 16882
rect 30770 16830 30782 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 34402 16830 34414 16882
rect 34466 16830 34478 16882
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 24894 16818 24946 16830
rect 30382 16818 30434 16830
rect 32510 16818 32562 16830
rect 38558 16818 38610 16830
rect 39006 16882 39058 16894
rect 39006 16818 39058 16830
rect 39342 16882 39394 16894
rect 39342 16818 39394 16830
rect 39678 16882 39730 16894
rect 39678 16818 39730 16830
rect 40462 16882 40514 16894
rect 40462 16818 40514 16830
rect 19070 16770 19122 16782
rect 19070 16706 19122 16718
rect 25678 16770 25730 16782
rect 37214 16770 37266 16782
rect 27794 16718 27806 16770
rect 27858 16718 27870 16770
rect 29922 16718 29934 16770
rect 29986 16718 29998 16770
rect 30818 16718 30830 16770
rect 30882 16718 30894 16770
rect 36530 16718 36542 16770
rect 36594 16718 36606 16770
rect 25678 16706 25730 16718
rect 37214 16706 37266 16718
rect 25902 16658 25954 16670
rect 25902 16594 25954 16606
rect 41806 16658 41858 16670
rect 41806 16594 41858 16606
rect 1344 16490 42560 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 42560 16490
rect 1344 16404 42560 16438
rect 33854 16322 33906 16334
rect 15362 16270 15374 16322
rect 15426 16319 15438 16322
rect 16258 16319 16270 16322
rect 15426 16273 16270 16319
rect 15426 16270 15438 16273
rect 16258 16270 16270 16273
rect 16322 16270 16334 16322
rect 20402 16270 20414 16322
rect 20466 16319 20478 16322
rect 20738 16319 20750 16322
rect 20466 16273 20750 16319
rect 20466 16270 20478 16273
rect 20738 16270 20750 16273
rect 20802 16270 20814 16322
rect 26786 16319 26798 16322
rect 26129 16273 26798 16319
rect 14366 16210 14418 16222
rect 14366 16146 14418 16158
rect 16270 16210 16322 16222
rect 16270 16146 16322 16158
rect 18734 16210 18786 16222
rect 18734 16146 18786 16158
rect 19182 16210 19234 16222
rect 19182 16146 19234 16158
rect 20414 16210 20466 16222
rect 20414 16146 20466 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 24670 16210 24722 16222
rect 24670 16146 24722 16158
rect 21982 16098 22034 16110
rect 21982 16034 22034 16046
rect 22318 16098 22370 16110
rect 22318 16034 22370 16046
rect 22990 16098 23042 16110
rect 22990 16034 23042 16046
rect 24110 16098 24162 16110
rect 24110 16034 24162 16046
rect 24334 16098 24386 16110
rect 24334 16034 24386 16046
rect 25454 16098 25506 16110
rect 25890 16046 25902 16098
rect 25954 16046 25966 16098
rect 25454 16034 25506 16046
rect 21646 15986 21698 15998
rect 21646 15922 21698 15934
rect 23102 15986 23154 15998
rect 23102 15922 23154 15934
rect 25230 15986 25282 15998
rect 26002 15934 26014 15986
rect 26066 15983 26078 15986
rect 26129 15983 26175 16273
rect 26786 16270 26798 16273
rect 26850 16270 26862 16322
rect 33854 16258 33906 16270
rect 39902 16322 39954 16334
rect 39902 16258 39954 16270
rect 26350 16210 26402 16222
rect 26350 16146 26402 16158
rect 27358 16210 27410 16222
rect 27358 16146 27410 16158
rect 28366 16210 28418 16222
rect 28366 16146 28418 16158
rect 30718 16210 30770 16222
rect 37662 16210 37714 16222
rect 39566 16210 39618 16222
rect 33170 16158 33182 16210
rect 33234 16158 33246 16210
rect 38770 16158 38782 16210
rect 38834 16158 38846 16210
rect 30718 16146 30770 16158
rect 37662 16146 37714 16158
rect 39566 16146 39618 16158
rect 27022 16098 27074 16110
rect 27022 16034 27074 16046
rect 27246 16098 27298 16110
rect 27246 16034 27298 16046
rect 27470 16098 27522 16110
rect 28254 16098 28306 16110
rect 30158 16098 30210 16110
rect 28018 16046 28030 16098
rect 28082 16046 28094 16098
rect 28690 16046 28702 16098
rect 28754 16046 28766 16098
rect 27470 16034 27522 16046
rect 28254 16034 28306 16046
rect 30158 16034 30210 16046
rect 31278 16098 31330 16110
rect 32846 16098 32898 16110
rect 31826 16046 31838 16098
rect 31890 16046 31902 16098
rect 31278 16034 31330 16046
rect 32846 16034 32898 16046
rect 33070 16098 33122 16110
rect 35310 16098 35362 16110
rect 33282 16046 33294 16098
rect 33346 16046 33358 16098
rect 33070 16034 33122 16046
rect 35310 16034 35362 16046
rect 35646 16098 35698 16110
rect 35646 16034 35698 16046
rect 35982 16098 36034 16110
rect 37438 16098 37490 16110
rect 36306 16046 36318 16098
rect 36370 16046 36382 16098
rect 35982 16034 36034 16046
rect 37438 16034 37490 16046
rect 39118 16098 39170 16110
rect 39118 16034 39170 16046
rect 41806 16098 41858 16110
rect 41806 16034 41858 16046
rect 26066 15937 26175 15983
rect 31502 15986 31554 15998
rect 26066 15934 26078 15937
rect 25230 15922 25282 15934
rect 31502 15922 31554 15934
rect 32622 15986 32674 15998
rect 32622 15922 32674 15934
rect 33966 15986 34018 15998
rect 33966 15922 34018 15934
rect 34638 15986 34690 15998
rect 34638 15922 34690 15934
rect 34750 15986 34802 15998
rect 34750 15922 34802 15934
rect 35422 15986 35474 15998
rect 35422 15922 35474 15934
rect 36542 15986 36594 15998
rect 36542 15922 36594 15934
rect 37998 15986 38050 15998
rect 37998 15922 38050 15934
rect 38782 15986 38834 15998
rect 38782 15922 38834 15934
rect 39790 15986 39842 15998
rect 39790 15922 39842 15934
rect 40574 15986 40626 15998
rect 40574 15922 40626 15934
rect 41694 15986 41746 15998
rect 41694 15922 41746 15934
rect 14926 15874 14978 15886
rect 14926 15810 14978 15822
rect 15374 15874 15426 15886
rect 15374 15810 15426 15822
rect 15710 15874 15762 15886
rect 15710 15810 15762 15822
rect 16718 15874 16770 15886
rect 16718 15810 16770 15822
rect 17166 15874 17218 15886
rect 17166 15810 17218 15822
rect 17614 15874 17666 15886
rect 17614 15810 17666 15822
rect 17950 15874 18002 15886
rect 17950 15810 18002 15822
rect 19742 15874 19794 15886
rect 19742 15810 19794 15822
rect 20862 15874 20914 15886
rect 20862 15810 20914 15822
rect 21982 15874 22034 15886
rect 21982 15810 22034 15822
rect 23326 15874 23378 15886
rect 23326 15810 23378 15822
rect 23438 15874 23490 15886
rect 23438 15810 23490 15822
rect 25566 15874 25618 15886
rect 25566 15810 25618 15822
rect 25678 15874 25730 15886
rect 25678 15810 25730 15822
rect 28478 15874 28530 15886
rect 28478 15810 28530 15822
rect 29486 15874 29538 15886
rect 29486 15810 29538 15822
rect 29598 15874 29650 15886
rect 29598 15810 29650 15822
rect 29822 15874 29874 15886
rect 29822 15810 29874 15822
rect 30606 15874 30658 15886
rect 30606 15810 30658 15822
rect 31390 15874 31442 15886
rect 31390 15810 31442 15822
rect 34414 15874 34466 15886
rect 34414 15810 34466 15822
rect 36654 15874 36706 15886
rect 36654 15810 36706 15822
rect 37774 15874 37826 15886
rect 37774 15810 37826 15822
rect 38558 15874 38610 15886
rect 38558 15810 38610 15822
rect 40462 15874 40514 15886
rect 40462 15810 40514 15822
rect 41022 15874 41074 15886
rect 41022 15810 41074 15822
rect 41470 15874 41522 15886
rect 42018 15822 42030 15874
rect 42082 15871 42094 15874
rect 42242 15871 42254 15874
rect 42082 15825 42254 15871
rect 42082 15822 42094 15825
rect 42242 15822 42254 15825
rect 42306 15822 42318 15874
rect 41470 15810 41522 15822
rect 1344 15706 42560 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 42560 15706
rect 1344 15620 42560 15654
rect 13358 15538 13410 15550
rect 13358 15474 13410 15486
rect 14590 15538 14642 15550
rect 14590 15474 14642 15486
rect 18286 15538 18338 15550
rect 18286 15474 18338 15486
rect 19966 15538 20018 15550
rect 19966 15474 20018 15486
rect 23886 15538 23938 15550
rect 23886 15474 23938 15486
rect 24110 15538 24162 15550
rect 24110 15474 24162 15486
rect 25902 15538 25954 15550
rect 25902 15474 25954 15486
rect 26910 15538 26962 15550
rect 26910 15474 26962 15486
rect 27134 15538 27186 15550
rect 27134 15474 27186 15486
rect 30382 15538 30434 15550
rect 30382 15474 30434 15486
rect 30606 15538 30658 15550
rect 30606 15474 30658 15486
rect 31502 15538 31554 15550
rect 31502 15474 31554 15486
rect 31614 15538 31666 15550
rect 31614 15474 31666 15486
rect 35646 15538 35698 15550
rect 35646 15474 35698 15486
rect 35870 15538 35922 15550
rect 35870 15474 35922 15486
rect 36430 15538 36482 15550
rect 36430 15474 36482 15486
rect 36654 15538 36706 15550
rect 36654 15474 36706 15486
rect 37214 15538 37266 15550
rect 37214 15474 37266 15486
rect 39790 15538 39842 15550
rect 39790 15474 39842 15486
rect 40574 15538 40626 15550
rect 40574 15474 40626 15486
rect 41806 15538 41858 15550
rect 41806 15474 41858 15486
rect 42030 15538 42082 15550
rect 42030 15474 42082 15486
rect 24222 15426 24274 15438
rect 21298 15374 21310 15426
rect 21362 15374 21374 15426
rect 24222 15362 24274 15374
rect 24670 15426 24722 15438
rect 24670 15362 24722 15374
rect 26238 15426 26290 15438
rect 26238 15362 26290 15374
rect 28702 15426 28754 15438
rect 28702 15362 28754 15374
rect 29486 15426 29538 15438
rect 29486 15362 29538 15374
rect 29934 15426 29986 15438
rect 29934 15362 29986 15374
rect 31726 15426 31778 15438
rect 31726 15362 31778 15374
rect 32398 15426 32450 15438
rect 32398 15362 32450 15374
rect 33742 15426 33794 15438
rect 33742 15362 33794 15374
rect 33854 15426 33906 15438
rect 33854 15362 33906 15374
rect 36318 15426 36370 15438
rect 36318 15362 36370 15374
rect 37102 15426 37154 15438
rect 37102 15362 37154 15374
rect 37438 15426 37490 15438
rect 37438 15362 37490 15374
rect 38334 15426 38386 15438
rect 38334 15362 38386 15374
rect 39454 15426 39506 15438
rect 39454 15362 39506 15374
rect 39566 15426 39618 15438
rect 39566 15362 39618 15374
rect 40350 15426 40402 15438
rect 40350 15362 40402 15374
rect 41694 15370 41746 15382
rect 25566 15314 25618 15326
rect 20626 15262 20638 15314
rect 20690 15262 20702 15314
rect 25566 15250 25618 15262
rect 26014 15314 26066 15326
rect 26014 15250 26066 15262
rect 26798 15314 26850 15326
rect 26798 15250 26850 15262
rect 27470 15314 27522 15326
rect 27470 15250 27522 15262
rect 28142 15314 28194 15326
rect 29374 15314 29426 15326
rect 30718 15314 30770 15326
rect 28466 15262 28478 15314
rect 28530 15262 28542 15314
rect 29698 15262 29710 15314
rect 29762 15262 29774 15314
rect 28142 15250 28194 15262
rect 29374 15250 29426 15262
rect 30718 15250 30770 15262
rect 32286 15314 32338 15326
rect 32286 15250 32338 15262
rect 33518 15314 33570 15326
rect 35534 15314 35586 15326
rect 34962 15262 34974 15314
rect 35026 15262 35038 15314
rect 33518 15250 33570 15262
rect 35534 15250 35586 15262
rect 38670 15314 38722 15326
rect 38670 15250 38722 15262
rect 38782 15314 38834 15326
rect 38782 15250 38834 15262
rect 38894 15314 38946 15326
rect 38894 15250 38946 15262
rect 40238 15314 40290 15326
rect 41694 15306 41746 15318
rect 40238 15250 40290 15262
rect 11678 15202 11730 15214
rect 11678 15138 11730 15150
rect 12574 15202 12626 15214
rect 12574 15138 12626 15150
rect 13022 15202 13074 15214
rect 13022 15138 13074 15150
rect 13918 15202 13970 15214
rect 13918 15138 13970 15150
rect 15262 15202 15314 15214
rect 15262 15138 15314 15150
rect 15822 15202 15874 15214
rect 15822 15138 15874 15150
rect 16494 15202 16546 15214
rect 16494 15138 16546 15150
rect 16942 15202 16994 15214
rect 16942 15138 16994 15150
rect 17838 15202 17890 15214
rect 17838 15138 17890 15150
rect 18846 15202 18898 15214
rect 18846 15138 18898 15150
rect 19182 15202 19234 15214
rect 28814 15202 28866 15214
rect 37774 15202 37826 15214
rect 23426 15150 23438 15202
rect 23490 15150 23502 15202
rect 34850 15150 34862 15202
rect 34914 15150 34926 15202
rect 19182 15138 19234 15150
rect 28814 15138 28866 15150
rect 37774 15138 37826 15150
rect 32398 15090 32450 15102
rect 24434 15038 24446 15090
rect 24498 15087 24510 15090
rect 25106 15087 25118 15090
rect 24498 15041 25118 15087
rect 24498 15038 24510 15041
rect 25106 15038 25118 15041
rect 25170 15038 25182 15090
rect 32398 15026 32450 15038
rect 1344 14922 42560 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 42560 14922
rect 1344 14836 42560 14870
rect 27246 14754 27298 14766
rect 11218 14702 11230 14754
rect 11282 14751 11294 14754
rect 11666 14751 11678 14754
rect 11282 14705 11678 14751
rect 11282 14702 11294 14705
rect 11666 14702 11678 14705
rect 11730 14702 11742 14754
rect 16930 14702 16942 14754
rect 16994 14751 17006 14754
rect 17266 14751 17278 14754
rect 16994 14705 17278 14751
rect 16994 14702 17006 14705
rect 17266 14702 17278 14705
rect 17330 14702 17342 14754
rect 27246 14690 27298 14702
rect 31278 14754 31330 14766
rect 31278 14690 31330 14702
rect 34190 14754 34242 14766
rect 34190 14690 34242 14702
rect 9662 14642 9714 14654
rect 9662 14578 9714 14590
rect 10110 14642 10162 14654
rect 10110 14578 10162 14590
rect 18622 14642 18674 14654
rect 25118 14642 25170 14654
rect 24546 14590 24558 14642
rect 24610 14590 24622 14642
rect 18622 14578 18674 14590
rect 25118 14578 25170 14590
rect 27918 14642 27970 14654
rect 34862 14642 34914 14654
rect 32722 14590 32734 14642
rect 32786 14590 32798 14642
rect 27918 14578 27970 14590
rect 34862 14578 34914 14590
rect 36206 14642 36258 14654
rect 36206 14578 36258 14590
rect 20078 14530 20130 14542
rect 27134 14530 27186 14542
rect 21746 14478 21758 14530
rect 21810 14478 21822 14530
rect 20078 14466 20130 14478
rect 27134 14466 27186 14478
rect 29598 14530 29650 14542
rect 29598 14466 29650 14478
rect 30270 14530 30322 14542
rect 30270 14466 30322 14478
rect 31390 14530 31442 14542
rect 31390 14466 31442 14478
rect 32398 14530 32450 14542
rect 32398 14466 32450 14478
rect 32622 14530 32674 14542
rect 33294 14530 33346 14542
rect 32834 14478 32846 14530
rect 32898 14478 32910 14530
rect 32622 14466 32674 14478
rect 33294 14466 33346 14478
rect 33630 14530 33682 14542
rect 33630 14466 33682 14478
rect 38782 14530 38834 14542
rect 38782 14466 38834 14478
rect 40350 14530 40402 14542
rect 40350 14466 40402 14478
rect 41806 14530 41858 14542
rect 41806 14466 41858 14478
rect 20190 14418 20242 14430
rect 26462 14418 26514 14430
rect 22418 14366 22430 14418
rect 22482 14366 22494 14418
rect 20190 14354 20242 14366
rect 26462 14354 26514 14366
rect 28814 14418 28866 14430
rect 28814 14354 28866 14366
rect 29710 14418 29762 14430
rect 29710 14354 29762 14366
rect 30606 14418 30658 14430
rect 30606 14354 30658 14366
rect 32174 14418 32226 14430
rect 32174 14354 32226 14366
rect 33518 14418 33570 14430
rect 33518 14354 33570 14366
rect 34302 14418 34354 14430
rect 34302 14354 34354 14366
rect 36094 14418 36146 14430
rect 36094 14354 36146 14366
rect 37662 14418 37714 14430
rect 37662 14354 37714 14366
rect 39118 14418 39170 14430
rect 39118 14354 39170 14366
rect 39566 14418 39618 14430
rect 40686 14418 40738 14430
rect 39890 14366 39902 14418
rect 39954 14366 39966 14418
rect 39566 14354 39618 14366
rect 40686 14354 40738 14366
rect 9214 14306 9266 14318
rect 9214 14242 9266 14254
rect 11118 14306 11170 14318
rect 11118 14242 11170 14254
rect 11566 14306 11618 14318
rect 11566 14242 11618 14254
rect 11902 14306 11954 14318
rect 11902 14242 11954 14254
rect 12462 14306 12514 14318
rect 12462 14242 12514 14254
rect 12910 14306 12962 14318
rect 12910 14242 12962 14254
rect 13582 14306 13634 14318
rect 13582 14242 13634 14254
rect 14142 14306 14194 14318
rect 14142 14242 14194 14254
rect 14478 14306 14530 14318
rect 14478 14242 14530 14254
rect 15038 14306 15090 14318
rect 15038 14242 15090 14254
rect 15598 14306 15650 14318
rect 15598 14242 15650 14254
rect 16046 14306 16098 14318
rect 16046 14242 16098 14254
rect 16494 14306 16546 14318
rect 16494 14242 16546 14254
rect 16942 14306 16994 14318
rect 16942 14242 16994 14254
rect 17390 14306 17442 14318
rect 17390 14242 17442 14254
rect 18174 14306 18226 14318
rect 18174 14242 18226 14254
rect 19070 14306 19122 14318
rect 19070 14242 19122 14254
rect 19630 14306 19682 14318
rect 19630 14242 19682 14254
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 20862 14306 20914 14318
rect 20862 14242 20914 14254
rect 25230 14306 25282 14318
rect 25230 14242 25282 14254
rect 25902 14306 25954 14318
rect 25902 14242 25954 14254
rect 26574 14306 26626 14318
rect 26574 14242 26626 14254
rect 27246 14306 27298 14318
rect 27246 14242 27298 14254
rect 28590 14306 28642 14318
rect 28590 14242 28642 14254
rect 28702 14306 28754 14318
rect 28702 14242 28754 14254
rect 29934 14306 29986 14318
rect 29934 14242 29986 14254
rect 30494 14306 30546 14318
rect 30494 14242 30546 14254
rect 31278 14306 31330 14318
rect 31278 14242 31330 14254
rect 34974 14306 35026 14318
rect 34974 14242 35026 14254
rect 35422 14306 35474 14318
rect 35422 14242 35474 14254
rect 36318 14306 36370 14318
rect 36318 14242 36370 14254
rect 36542 14306 36594 14318
rect 36542 14242 36594 14254
rect 37550 14306 37602 14318
rect 37550 14242 37602 14254
rect 38110 14306 38162 14318
rect 38110 14242 38162 14254
rect 38894 14306 38946 14318
rect 38894 14242 38946 14254
rect 40574 14306 40626 14318
rect 40574 14242 40626 14254
rect 41470 14306 41522 14318
rect 41470 14242 41522 14254
rect 41694 14306 41746 14318
rect 41694 14242 41746 14254
rect 1344 14138 42560 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 42560 14138
rect 1344 14052 42560 14086
rect 15150 13970 15202 13982
rect 15150 13906 15202 13918
rect 15598 13970 15650 13982
rect 15598 13906 15650 13918
rect 16606 13970 16658 13982
rect 16606 13906 16658 13918
rect 16942 13970 16994 13982
rect 16942 13906 16994 13918
rect 24110 13970 24162 13982
rect 24110 13906 24162 13918
rect 27022 13970 27074 13982
rect 27022 13906 27074 13918
rect 32734 13970 32786 13982
rect 32734 13906 32786 13918
rect 33854 13970 33906 13982
rect 33854 13906 33906 13918
rect 34862 13970 34914 13982
rect 34862 13906 34914 13918
rect 36206 13970 36258 13982
rect 39454 13970 39506 13982
rect 36642 13918 36654 13970
rect 36706 13918 36718 13970
rect 36206 13906 36258 13918
rect 39454 13906 39506 13918
rect 39566 13970 39618 13982
rect 39566 13906 39618 13918
rect 40014 13970 40066 13982
rect 40014 13906 40066 13918
rect 41694 13970 41746 13982
rect 41694 13906 41746 13918
rect 14254 13858 14306 13870
rect 14254 13794 14306 13806
rect 21310 13858 21362 13870
rect 21310 13794 21362 13806
rect 21534 13858 21586 13870
rect 21534 13794 21586 13806
rect 21646 13858 21698 13870
rect 21646 13794 21698 13806
rect 22766 13858 22818 13870
rect 22766 13794 22818 13806
rect 24782 13858 24834 13870
rect 24782 13794 24834 13806
rect 28478 13858 28530 13870
rect 28478 13794 28530 13806
rect 32510 13858 32562 13870
rect 32510 13794 32562 13806
rect 32846 13858 32898 13870
rect 32846 13794 32898 13806
rect 33630 13858 33682 13870
rect 33630 13794 33682 13806
rect 35982 13858 36034 13870
rect 35982 13794 36034 13806
rect 37214 13858 37266 13870
rect 37214 13794 37266 13806
rect 38334 13858 38386 13870
rect 38334 13794 38386 13806
rect 40686 13858 40738 13870
rect 40686 13794 40738 13806
rect 13358 13746 13410 13758
rect 22878 13746 22930 13758
rect 17938 13694 17950 13746
rect 18002 13694 18014 13746
rect 21970 13694 21982 13746
rect 22034 13694 22046 13746
rect 13358 13682 13410 13694
rect 22878 13682 22930 13694
rect 24894 13746 24946 13758
rect 24894 13682 24946 13694
rect 25678 13746 25730 13758
rect 25678 13682 25730 13694
rect 25902 13746 25954 13758
rect 25902 13682 25954 13694
rect 26350 13746 26402 13758
rect 26350 13682 26402 13694
rect 26798 13746 26850 13758
rect 26798 13682 26850 13694
rect 26910 13746 26962 13758
rect 34078 13746 34130 13758
rect 35870 13746 35922 13758
rect 27346 13694 27358 13746
rect 27410 13694 27422 13746
rect 28018 13694 28030 13746
rect 28082 13694 28094 13746
rect 29250 13694 29262 13746
rect 29314 13694 29326 13746
rect 34290 13694 34302 13746
rect 34354 13694 34366 13746
rect 26910 13682 26962 13694
rect 34078 13682 34130 13694
rect 35870 13682 35922 13694
rect 38894 13746 38946 13758
rect 38894 13682 38946 13694
rect 39342 13746 39394 13758
rect 39342 13682 39394 13694
rect 40574 13746 40626 13758
rect 40574 13682 40626 13694
rect 40910 13746 40962 13758
rect 40910 13682 40962 13694
rect 41582 13746 41634 13758
rect 41582 13682 41634 13694
rect 6750 13634 6802 13646
rect 6750 13570 6802 13582
rect 7198 13634 7250 13646
rect 7198 13570 7250 13582
rect 7646 13634 7698 13646
rect 7646 13570 7698 13582
rect 8094 13634 8146 13646
rect 8094 13570 8146 13582
rect 8654 13634 8706 13646
rect 8654 13570 8706 13582
rect 8990 13634 9042 13646
rect 8990 13570 9042 13582
rect 9886 13634 9938 13646
rect 9886 13570 9938 13582
rect 10334 13634 10386 13646
rect 10334 13570 10386 13582
rect 11118 13634 11170 13646
rect 11118 13570 11170 13582
rect 11678 13634 11730 13646
rect 11678 13570 11730 13582
rect 12014 13634 12066 13646
rect 12014 13570 12066 13582
rect 12574 13634 12626 13646
rect 12574 13570 12626 13582
rect 12910 13634 12962 13646
rect 12910 13570 12962 13582
rect 13918 13634 13970 13646
rect 13918 13570 13970 13582
rect 14702 13634 14754 13646
rect 14702 13570 14754 13582
rect 16046 13634 16098 13646
rect 23550 13634 23602 13646
rect 18610 13582 18622 13634
rect 18674 13582 18686 13634
rect 20738 13582 20750 13634
rect 20802 13582 20814 13634
rect 22082 13582 22094 13634
rect 22146 13582 22158 13634
rect 16046 13570 16098 13582
rect 23550 13570 23602 13582
rect 25790 13634 25842 13646
rect 33966 13634 34018 13646
rect 29922 13582 29934 13634
rect 29986 13582 29998 13634
rect 32050 13582 32062 13634
rect 32114 13582 32126 13634
rect 25790 13570 25842 13582
rect 33966 13570 34018 13582
rect 34974 13634 35026 13646
rect 38434 13582 38446 13634
rect 38498 13582 38510 13634
rect 34974 13570 35026 13582
rect 22766 13522 22818 13534
rect 6738 13470 6750 13522
rect 6802 13519 6814 13522
rect 7410 13519 7422 13522
rect 6802 13473 7422 13519
rect 6802 13470 6814 13473
rect 7410 13470 7422 13473
rect 7474 13470 7486 13522
rect 7634 13470 7646 13522
rect 7698 13519 7710 13522
rect 8866 13519 8878 13522
rect 7698 13473 8878 13519
rect 7698 13470 7710 13473
rect 8866 13470 8878 13473
rect 8930 13519 8942 13522
rect 9202 13519 9214 13522
rect 8930 13473 9214 13519
rect 8930 13470 8942 13473
rect 9202 13470 9214 13473
rect 9266 13470 9278 13522
rect 12562 13470 12574 13522
rect 12626 13519 12638 13522
rect 13234 13519 13246 13522
rect 12626 13473 13246 13519
rect 12626 13470 12638 13473
rect 13234 13470 13246 13473
rect 13298 13470 13310 13522
rect 13570 13470 13582 13522
rect 13634 13519 13646 13522
rect 14130 13519 14142 13522
rect 13634 13473 14142 13519
rect 13634 13470 13646 13473
rect 14130 13470 14142 13473
rect 14194 13470 14206 13522
rect 16146 13470 16158 13522
rect 16210 13519 16222 13522
rect 16594 13519 16606 13522
rect 16210 13473 16606 13519
rect 16210 13470 16222 13473
rect 16594 13470 16606 13473
rect 16658 13470 16670 13522
rect 22766 13458 22818 13470
rect 24782 13522 24834 13534
rect 24782 13458 24834 13470
rect 36990 13522 37042 13534
rect 36990 13458 37042 13470
rect 38110 13522 38162 13534
rect 38110 13458 38162 13470
rect 41694 13522 41746 13534
rect 41694 13458 41746 13470
rect 1344 13354 42560 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 42560 13354
rect 1344 13268 42560 13302
rect 27806 13186 27858 13198
rect 27806 13122 27858 13134
rect 36654 13186 36706 13198
rect 36654 13122 36706 13134
rect 6414 13074 6466 13086
rect 12686 13074 12738 13086
rect 22990 13074 23042 13086
rect 29710 13074 29762 13086
rect 37774 13074 37826 13086
rect 7186 13022 7198 13074
rect 7250 13022 7262 13074
rect 20402 13022 20414 13074
rect 20466 13022 20478 13074
rect 27122 13022 27134 13074
rect 27186 13022 27198 13074
rect 33058 13022 33070 13074
rect 33122 13022 33134 13074
rect 35186 13022 35198 13074
rect 35250 13022 35262 13074
rect 6414 13010 6466 13022
rect 12686 13010 12738 13022
rect 22990 13010 23042 13022
rect 29710 13010 29762 13022
rect 37774 13010 37826 13022
rect 12126 12962 12178 12974
rect 10098 12910 10110 12962
rect 10162 12910 10174 12962
rect 12126 12898 12178 12910
rect 13694 12962 13746 12974
rect 13694 12898 13746 12910
rect 19070 12962 19122 12974
rect 19070 12898 19122 12910
rect 19742 12962 19794 12974
rect 29486 12962 29538 12974
rect 20738 12910 20750 12962
rect 20802 12910 20814 12962
rect 23426 12910 23438 12962
rect 23490 12910 23502 12962
rect 24210 12910 24222 12962
rect 24274 12910 24286 12962
rect 19742 12898 19794 12910
rect 29486 12898 29538 12910
rect 30158 12962 30210 12974
rect 30158 12898 30210 12910
rect 31054 12962 31106 12974
rect 35758 12962 35810 12974
rect 32386 12910 32398 12962
rect 32450 12910 32462 12962
rect 31054 12898 31106 12910
rect 35758 12898 35810 12910
rect 38222 12962 38274 12974
rect 38222 12898 38274 12910
rect 38670 12962 38722 12974
rect 38670 12898 38722 12910
rect 39342 12962 39394 12974
rect 39342 12898 39394 12910
rect 39678 12962 39730 12974
rect 39678 12898 39730 12910
rect 40014 12962 40066 12974
rect 40014 12898 40066 12910
rect 40574 12962 40626 12974
rect 40574 12898 40626 12910
rect 41470 12962 41522 12974
rect 41470 12898 41522 12910
rect 41806 12962 41858 12974
rect 41806 12898 41858 12910
rect 10782 12850 10834 12862
rect 9314 12798 9326 12850
rect 9378 12798 9390 12850
rect 10782 12786 10834 12798
rect 12014 12850 12066 12862
rect 12014 12786 12066 12798
rect 12798 12850 12850 12862
rect 14478 12850 14530 12862
rect 12898 12798 12910 12850
rect 12962 12847 12974 12850
rect 13122 12847 13134 12850
rect 12962 12801 13134 12847
rect 12962 12798 12974 12801
rect 13122 12798 13134 12801
rect 13186 12798 13198 12850
rect 12798 12786 12850 12798
rect 14478 12786 14530 12798
rect 17278 12850 17330 12862
rect 17278 12786 17330 12798
rect 17838 12850 17890 12862
rect 17838 12786 17890 12798
rect 18510 12850 18562 12862
rect 18510 12786 18562 12798
rect 21982 12850 22034 12862
rect 27694 12850 27746 12862
rect 24994 12798 25006 12850
rect 25058 12798 25070 12850
rect 21982 12786 22034 12798
rect 27694 12786 27746 12798
rect 28366 12850 28418 12862
rect 28366 12786 28418 12798
rect 29934 12850 29986 12862
rect 29934 12786 29986 12798
rect 30718 12850 30770 12862
rect 30718 12786 30770 12798
rect 30830 12850 30882 12862
rect 30830 12786 30882 12798
rect 31502 12850 31554 12862
rect 31502 12786 31554 12798
rect 31614 12850 31666 12862
rect 31614 12786 31666 12798
rect 35870 12850 35922 12862
rect 35870 12786 35922 12798
rect 36094 12850 36146 12862
rect 36094 12786 36146 12798
rect 36654 12850 36706 12862
rect 36654 12786 36706 12798
rect 36766 12850 36818 12862
rect 36766 12786 36818 12798
rect 37662 12850 37714 12862
rect 37662 12786 37714 12798
rect 37998 12850 38050 12862
rect 37998 12786 38050 12798
rect 39006 12850 39058 12862
rect 39006 12786 39058 12798
rect 39902 12850 39954 12862
rect 39902 12786 39954 12798
rect 5966 12738 6018 12750
rect 5966 12674 6018 12686
rect 10670 12738 10722 12750
rect 10670 12674 10722 12686
rect 11454 12738 11506 12750
rect 11454 12674 11506 12686
rect 13806 12738 13858 12750
rect 13806 12674 13858 12686
rect 14030 12738 14082 12750
rect 14030 12674 14082 12686
rect 14590 12738 14642 12750
rect 14590 12674 14642 12686
rect 15486 12738 15538 12750
rect 15486 12674 15538 12686
rect 15934 12738 15986 12750
rect 15934 12674 15986 12686
rect 16270 12738 16322 12750
rect 16270 12674 16322 12686
rect 16830 12738 16882 12750
rect 16830 12674 16882 12686
rect 17726 12738 17778 12750
rect 17726 12674 17778 12686
rect 18398 12738 18450 12750
rect 18398 12674 18450 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 22094 12738 22146 12750
rect 22094 12674 22146 12686
rect 22878 12738 22930 12750
rect 22878 12674 22930 12686
rect 23102 12738 23154 12750
rect 23102 12674 23154 12686
rect 27918 12738 27970 12750
rect 27918 12674 27970 12686
rect 28142 12738 28194 12750
rect 28142 12674 28194 12686
rect 28814 12738 28866 12750
rect 28814 12674 28866 12686
rect 31838 12738 31890 12750
rect 31838 12674 31890 12686
rect 38782 12738 38834 12750
rect 38782 12674 38834 12686
rect 40686 12738 40738 12750
rect 40686 12674 40738 12686
rect 40910 12738 40962 12750
rect 40910 12674 40962 12686
rect 41694 12738 41746 12750
rect 41694 12674 41746 12686
rect 1344 12570 42560 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 42560 12570
rect 1344 12484 42560 12518
rect 12798 12402 12850 12414
rect 12798 12338 12850 12350
rect 15150 12402 15202 12414
rect 15150 12338 15202 12350
rect 15822 12402 15874 12414
rect 15822 12338 15874 12350
rect 16382 12402 16434 12414
rect 30606 12402 30658 12414
rect 29474 12350 29486 12402
rect 29538 12350 29550 12402
rect 16382 12338 16434 12350
rect 30606 12338 30658 12350
rect 32846 12402 32898 12414
rect 32846 12338 32898 12350
rect 33742 12402 33794 12414
rect 33742 12338 33794 12350
rect 35534 12402 35586 12414
rect 35534 12338 35586 12350
rect 36430 12402 36482 12414
rect 36430 12338 36482 12350
rect 36654 12402 36706 12414
rect 36654 12338 36706 12350
rect 37438 12402 37490 12414
rect 37438 12338 37490 12350
rect 38222 12402 38274 12414
rect 38222 12338 38274 12350
rect 38446 12402 38498 12414
rect 38446 12338 38498 12350
rect 39678 12402 39730 12414
rect 39678 12338 39730 12350
rect 41694 12402 41746 12414
rect 41694 12338 41746 12350
rect 9886 12290 9938 12302
rect 9886 12226 9938 12238
rect 11902 12290 11954 12302
rect 11902 12226 11954 12238
rect 13470 12290 13522 12302
rect 13470 12226 13522 12238
rect 13582 12290 13634 12302
rect 13582 12226 13634 12238
rect 14254 12290 14306 12302
rect 14254 12226 14306 12238
rect 14366 12290 14418 12302
rect 14366 12226 14418 12238
rect 15038 12290 15090 12302
rect 15038 12226 15090 12238
rect 18846 12290 18898 12302
rect 18846 12226 18898 12238
rect 18958 12290 19010 12302
rect 18958 12226 19010 12238
rect 25790 12290 25842 12302
rect 25790 12226 25842 12238
rect 25902 12290 25954 12302
rect 25902 12226 25954 12238
rect 27582 12290 27634 12302
rect 27582 12226 27634 12238
rect 28254 12290 28306 12302
rect 28254 12226 28306 12238
rect 28926 12290 28978 12302
rect 28926 12226 28978 12238
rect 29822 12290 29874 12302
rect 29822 12226 29874 12238
rect 33630 12290 33682 12302
rect 34526 12290 34578 12302
rect 34290 12238 34302 12290
rect 34354 12238 34366 12290
rect 33630 12226 33682 12238
rect 34526 12226 34578 12238
rect 35086 12290 35138 12302
rect 35086 12226 35138 12238
rect 36766 12290 36818 12302
rect 36766 12226 36818 12238
rect 37326 12290 37378 12302
rect 37326 12226 37378 12238
rect 38670 12290 38722 12302
rect 38670 12226 38722 12238
rect 39454 12290 39506 12302
rect 39454 12226 39506 12238
rect 40462 12290 40514 12302
rect 40462 12226 40514 12238
rect 40574 12290 40626 12302
rect 40574 12226 40626 12238
rect 41806 12290 41858 12302
rect 41806 12226 41858 12238
rect 10222 12178 10274 12190
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 10222 12114 10274 12126
rect 11006 12178 11058 12190
rect 11006 12114 11058 12126
rect 12574 12178 12626 12190
rect 12574 12114 12626 12126
rect 12910 12178 12962 12190
rect 12910 12114 12962 12126
rect 14590 12178 14642 12190
rect 14590 12114 14642 12126
rect 15374 12178 15426 12190
rect 15374 12114 15426 12126
rect 19182 12178 19234 12190
rect 25566 12178 25618 12190
rect 23650 12126 23662 12178
rect 23714 12126 23726 12178
rect 19182 12114 19234 12126
rect 25566 12114 25618 12126
rect 26910 12178 26962 12190
rect 26910 12114 26962 12126
rect 27358 12178 27410 12190
rect 27358 12114 27410 12126
rect 28366 12178 28418 12190
rect 28366 12114 28418 12126
rect 29150 12178 29202 12190
rect 30942 12178 30994 12190
rect 29586 12126 29598 12178
rect 29650 12126 29662 12178
rect 30482 12126 30494 12178
rect 30546 12126 30558 12178
rect 29150 12114 29202 12126
rect 30942 12114 30994 12126
rect 31838 12178 31890 12190
rect 31838 12114 31890 12126
rect 33854 12178 33906 12190
rect 33854 12114 33906 12126
rect 35310 12178 35362 12190
rect 36094 12178 36146 12190
rect 35746 12126 35758 12178
rect 35810 12126 35822 12178
rect 35310 12114 35362 12126
rect 36094 12114 36146 12126
rect 4734 12066 4786 12078
rect 4734 12002 4786 12014
rect 5070 12066 5122 12078
rect 5070 12002 5122 12014
rect 5630 12066 5682 12078
rect 11118 12066 11170 12078
rect 6850 12014 6862 12066
rect 6914 12014 6926 12066
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 5630 12002 5682 12014
rect 11118 12002 11170 12014
rect 12126 12066 12178 12078
rect 12126 12002 12178 12014
rect 16830 12066 16882 12078
rect 16830 12002 16882 12014
rect 17614 12066 17666 12078
rect 17614 12002 17666 12014
rect 18286 12066 18338 12078
rect 30718 12066 30770 12078
rect 21746 12014 21758 12066
rect 21810 12014 21822 12066
rect 32274 12014 32286 12066
rect 32338 12014 32350 12066
rect 39778 12014 39790 12066
rect 39842 12014 39854 12066
rect 18286 12002 18338 12014
rect 30718 12002 30770 12014
rect 9998 11954 10050 11966
rect 9998 11890 10050 11902
rect 10334 11954 10386 11966
rect 10334 11890 10386 11902
rect 11790 11954 11842 11966
rect 11790 11890 11842 11902
rect 13582 11954 13634 11966
rect 13582 11890 13634 11902
rect 16942 11954 16994 11966
rect 18174 11954 18226 11966
rect 17602 11902 17614 11954
rect 17666 11951 17678 11954
rect 17938 11951 17950 11954
rect 17666 11905 17950 11951
rect 17666 11902 17678 11905
rect 17938 11902 17950 11905
rect 18002 11902 18014 11954
rect 16942 11890 16994 11902
rect 18174 11890 18226 11902
rect 26462 11954 26514 11966
rect 26462 11890 26514 11902
rect 27134 11954 27186 11966
rect 27134 11890 27186 11902
rect 28254 11954 28306 11966
rect 28254 11890 28306 11902
rect 29374 11954 29426 11966
rect 29374 11890 29426 11902
rect 31166 11954 31218 11966
rect 31166 11890 31218 11902
rect 34078 11954 34130 11966
rect 34078 11890 34130 11902
rect 35534 11954 35586 11966
rect 35534 11890 35586 11902
rect 37438 11954 37490 11966
rect 37438 11890 37490 11902
rect 38110 11954 38162 11966
rect 38110 11890 38162 11902
rect 40462 11954 40514 11966
rect 40462 11890 40514 11902
rect 41694 11954 41746 11966
rect 41694 11890 41746 11902
rect 1344 11786 42560 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 42560 11786
rect 1344 11700 42560 11734
rect 9662 11618 9714 11630
rect 9662 11554 9714 11566
rect 11006 11618 11058 11630
rect 11006 11554 11058 11566
rect 12798 11618 12850 11630
rect 12798 11554 12850 11566
rect 14814 11618 14866 11630
rect 14814 11554 14866 11566
rect 22542 11618 22594 11630
rect 22542 11554 22594 11566
rect 40462 11618 40514 11630
rect 40462 11554 40514 11566
rect 41918 11618 41970 11630
rect 41918 11554 41970 11566
rect 6862 11506 6914 11518
rect 11790 11506 11842 11518
rect 28702 11506 28754 11518
rect 36766 11506 36818 11518
rect 42030 11506 42082 11518
rect 9874 11454 9886 11506
rect 9938 11454 9950 11506
rect 13906 11454 13918 11506
rect 13970 11454 13982 11506
rect 19394 11454 19406 11506
rect 19458 11454 19470 11506
rect 24210 11454 24222 11506
rect 24274 11454 24286 11506
rect 32162 11454 32174 11506
rect 32226 11454 32238 11506
rect 39442 11454 39454 11506
rect 39506 11454 39518 11506
rect 6862 11442 6914 11454
rect 11790 11442 11842 11454
rect 28702 11442 28754 11454
rect 36766 11442 36818 11454
rect 42030 11442 42082 11454
rect 7758 11394 7810 11406
rect 7074 11342 7086 11394
rect 7138 11342 7150 11394
rect 7758 11330 7810 11342
rect 10894 11394 10946 11406
rect 10894 11330 10946 11342
rect 15934 11394 15986 11406
rect 19966 11394 20018 11406
rect 16594 11342 16606 11394
rect 16658 11342 16670 11394
rect 15934 11330 15986 11342
rect 19966 11330 20018 11342
rect 20190 11394 20242 11406
rect 20190 11330 20242 11342
rect 21870 11394 21922 11406
rect 32846 11394 32898 11406
rect 26898 11342 26910 11394
rect 26962 11342 26974 11394
rect 30146 11342 30158 11394
rect 30210 11342 30222 11394
rect 21870 11330 21922 11342
rect 32846 11330 32898 11342
rect 34638 11394 34690 11406
rect 34638 11330 34690 11342
rect 34862 11394 34914 11406
rect 34862 11330 34914 11342
rect 35086 11394 35138 11406
rect 37774 11394 37826 11406
rect 36082 11342 36094 11394
rect 36146 11342 36158 11394
rect 35086 11330 35138 11342
rect 37774 11330 37826 11342
rect 38222 11394 38274 11406
rect 38222 11330 38274 11342
rect 39790 11394 39842 11406
rect 39790 11330 39842 11342
rect 41358 11394 41410 11406
rect 41358 11330 41410 11342
rect 6078 11282 6130 11294
rect 6078 11218 6130 11230
rect 6750 11282 6802 11294
rect 6750 11218 6802 11230
rect 8094 11282 8146 11294
rect 8094 11218 8146 11230
rect 8654 11282 8706 11294
rect 8654 11218 8706 11230
rect 8990 11282 9042 11294
rect 8990 11218 9042 11230
rect 11678 11282 11730 11294
rect 11678 11218 11730 11230
rect 12126 11282 12178 11294
rect 12126 11218 12178 11230
rect 12910 11282 12962 11294
rect 12910 11218 12962 11230
rect 14142 11282 14194 11294
rect 14142 11218 14194 11230
rect 14702 11282 14754 11294
rect 31390 11282 31442 11294
rect 17266 11230 17278 11282
rect 17330 11230 17342 11282
rect 29586 11230 29598 11282
rect 29650 11230 29662 11282
rect 14702 11218 14754 11230
rect 31390 11218 31442 11230
rect 31950 11282 32002 11294
rect 31950 11218 32002 11230
rect 32958 11282 33010 11294
rect 32958 11218 33010 11230
rect 34190 11282 34242 11294
rect 37662 11282 37714 11294
rect 34402 11230 34414 11282
rect 34466 11230 34478 11282
rect 34190 11218 34242 11230
rect 37662 11218 37714 11230
rect 38446 11282 38498 11294
rect 38446 11218 38498 11230
rect 38558 11282 38610 11294
rect 38558 11218 38610 11230
rect 40462 11282 40514 11294
rect 40462 11218 40514 11230
rect 40574 11282 40626 11294
rect 40574 11218 40626 11230
rect 41246 11282 41298 11294
rect 41246 11218 41298 11230
rect 3614 11170 3666 11182
rect 3614 11106 3666 11118
rect 4062 11170 4114 11182
rect 4062 11106 4114 11118
rect 4510 11170 4562 11182
rect 4510 11106 4562 11118
rect 4958 11170 5010 11182
rect 4958 11106 5010 11118
rect 6190 11170 6242 11182
rect 6190 11106 6242 11118
rect 7646 11170 7698 11182
rect 7646 11106 7698 11118
rect 7870 11170 7922 11182
rect 7870 11106 7922 11118
rect 8878 11170 8930 11182
rect 8878 11106 8930 11118
rect 9886 11170 9938 11182
rect 9886 11106 9938 11118
rect 11006 11170 11058 11182
rect 11006 11106 11058 11118
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 13918 11170 13970 11182
rect 13918 11106 13970 11118
rect 15374 11170 15426 11182
rect 22206 11170 22258 11182
rect 20514 11118 20526 11170
rect 20578 11118 20590 11170
rect 15374 11106 15426 11118
rect 22206 11106 22258 11118
rect 22430 11170 22482 11182
rect 30830 11170 30882 11182
rect 30034 11118 30046 11170
rect 30098 11118 30110 11170
rect 22430 11106 22482 11118
rect 30830 11106 30882 11118
rect 33182 11170 33234 11182
rect 33182 11106 33234 11118
rect 33518 11170 33570 11182
rect 36094 11170 36146 11182
rect 34514 11118 34526 11170
rect 34578 11118 34590 11170
rect 33518 11106 33570 11118
rect 36094 11106 36146 11118
rect 37438 11170 37490 11182
rect 37438 11106 37490 11118
rect 39566 11170 39618 11182
rect 39566 11106 39618 11118
rect 41022 11170 41074 11182
rect 41022 11106 41074 11118
rect 1344 11002 42560 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 42560 11002
rect 1344 10916 42560 10950
rect 2718 10834 2770 10846
rect 2718 10770 2770 10782
rect 4398 10834 4450 10846
rect 4398 10770 4450 10782
rect 8430 10834 8482 10846
rect 8430 10770 8482 10782
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 23550 10834 23602 10846
rect 23550 10770 23602 10782
rect 24334 10834 24386 10846
rect 29822 10834 29874 10846
rect 26674 10782 26686 10834
rect 26738 10782 26750 10834
rect 24334 10770 24386 10782
rect 29822 10770 29874 10782
rect 30494 10834 30546 10846
rect 30494 10770 30546 10782
rect 31166 10834 31218 10846
rect 31166 10770 31218 10782
rect 32286 10834 32338 10846
rect 32286 10770 32338 10782
rect 32622 10834 32674 10846
rect 32622 10770 32674 10782
rect 34302 10834 34354 10846
rect 34302 10770 34354 10782
rect 35982 10834 36034 10846
rect 35982 10770 36034 10782
rect 38334 10834 38386 10846
rect 38334 10770 38386 10782
rect 39230 10834 39282 10846
rect 39230 10770 39282 10782
rect 40238 10834 40290 10846
rect 40238 10770 40290 10782
rect 41694 10834 41746 10846
rect 41694 10770 41746 10782
rect 6302 10722 6354 10734
rect 6302 10658 6354 10670
rect 7646 10722 7698 10734
rect 7646 10658 7698 10670
rect 9886 10722 9938 10734
rect 9886 10658 9938 10670
rect 9998 10722 10050 10734
rect 14702 10722 14754 10734
rect 13010 10670 13022 10722
rect 13074 10670 13086 10722
rect 9998 10658 10050 10670
rect 14702 10658 14754 10670
rect 16942 10722 16994 10734
rect 16942 10658 16994 10670
rect 18174 10722 18226 10734
rect 18174 10658 18226 10670
rect 18846 10722 18898 10734
rect 18846 10658 18898 10670
rect 19070 10722 19122 10734
rect 19070 10658 19122 10670
rect 23438 10722 23490 10734
rect 23438 10658 23490 10670
rect 24558 10722 24610 10734
rect 27918 10722 27970 10734
rect 25890 10670 25902 10722
rect 25954 10670 25966 10722
rect 26562 10670 26574 10722
rect 26626 10670 26638 10722
rect 24558 10658 24610 10670
rect 27918 10658 27970 10670
rect 28366 10722 28418 10734
rect 28366 10658 28418 10670
rect 28590 10722 28642 10734
rect 28590 10658 28642 10670
rect 31390 10722 31442 10734
rect 31390 10658 31442 10670
rect 32062 10722 32114 10734
rect 32062 10658 32114 10670
rect 33742 10722 33794 10734
rect 33742 10658 33794 10670
rect 35870 10722 35922 10734
rect 35870 10658 35922 10670
rect 39342 10722 39394 10734
rect 39342 10658 39394 10670
rect 40350 10722 40402 10734
rect 40350 10658 40402 10670
rect 41806 10722 41858 10734
rect 41806 10658 41858 10670
rect 6862 10610 6914 10622
rect 6862 10546 6914 10558
rect 8318 10610 8370 10622
rect 14366 10610 14418 10622
rect 13794 10558 13806 10610
rect 13858 10558 13870 10610
rect 8318 10546 8370 10558
rect 14366 10546 14418 10558
rect 16830 10610 16882 10622
rect 24222 10610 24274 10622
rect 28702 10610 28754 10622
rect 31502 10610 31554 10622
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 24770 10558 24782 10610
rect 24834 10558 24846 10610
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 27458 10558 27470 10610
rect 27522 10558 27534 10610
rect 30594 10558 30606 10610
rect 30658 10558 30670 10610
rect 16830 10546 16882 10558
rect 24222 10546 24274 10558
rect 28702 10546 28754 10558
rect 31502 10546 31554 10558
rect 32510 10610 32562 10622
rect 32510 10546 32562 10558
rect 33630 10610 33682 10622
rect 33630 10546 33682 10558
rect 34414 10610 34466 10622
rect 34414 10546 34466 10558
rect 34974 10610 35026 10622
rect 34974 10546 35026 10558
rect 35422 10610 35474 10622
rect 35422 10546 35474 10558
rect 37438 10610 37490 10622
rect 37438 10546 37490 10558
rect 37662 10610 37714 10622
rect 37662 10546 37714 10558
rect 38110 10610 38162 10622
rect 38110 10546 38162 10558
rect 38446 10610 38498 10622
rect 38446 10546 38498 10558
rect 38670 10610 38722 10622
rect 39554 10558 39566 10610
rect 39618 10558 39630 10610
rect 39778 10558 39790 10610
rect 39842 10558 39854 10610
rect 40562 10558 40574 10610
rect 40626 10558 40638 10610
rect 40786 10558 40798 10610
rect 40850 10558 40862 10610
rect 38670 10546 38722 10558
rect 3166 10498 3218 10510
rect 3166 10434 3218 10446
rect 3502 10498 3554 10510
rect 3502 10434 3554 10446
rect 4062 10498 4114 10510
rect 4062 10434 4114 10446
rect 4846 10498 4898 10510
rect 4846 10434 4898 10446
rect 5294 10498 5346 10510
rect 5294 10434 5346 10446
rect 5742 10498 5794 10510
rect 5742 10434 5794 10446
rect 7534 10498 7586 10510
rect 7534 10434 7586 10446
rect 8990 10498 9042 10510
rect 15486 10498 15538 10510
rect 29262 10498 29314 10510
rect 34638 10498 34690 10510
rect 10882 10446 10894 10498
rect 10946 10446 10958 10498
rect 15810 10446 15822 10498
rect 15874 10446 15886 10498
rect 17938 10446 17950 10498
rect 18002 10446 18014 10498
rect 20738 10446 20750 10498
rect 20802 10446 20814 10498
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 32610 10446 32622 10498
rect 32674 10446 32686 10498
rect 8990 10434 9042 10446
rect 15486 10434 15538 10446
rect 29262 10434 29314 10446
rect 34638 10434 34690 10446
rect 36542 10498 36594 10510
rect 36542 10434 36594 10446
rect 37102 10498 37154 10510
rect 37102 10434 37154 10446
rect 6750 10386 6802 10398
rect 6750 10322 6802 10334
rect 7422 10386 7474 10398
rect 7422 10322 7474 10334
rect 8430 10386 8482 10398
rect 8430 10322 8482 10334
rect 9886 10386 9938 10398
rect 9886 10322 9938 10334
rect 16494 10386 16546 10398
rect 16494 10322 16546 10334
rect 16606 10386 16658 10398
rect 16606 10322 16658 10334
rect 18734 10386 18786 10398
rect 18734 10322 18786 10334
rect 33742 10386 33794 10398
rect 33742 10322 33794 10334
rect 34862 10386 34914 10398
rect 34862 10322 34914 10334
rect 35982 10386 36034 10398
rect 35982 10322 36034 10334
rect 41694 10386 41746 10398
rect 41694 10322 41746 10334
rect 1344 10218 42560 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 42560 10218
rect 1344 10132 42560 10166
rect 10446 10050 10498 10062
rect 2370 9998 2382 10050
rect 2434 10047 2446 10050
rect 3154 10047 3166 10050
rect 2434 10001 3166 10047
rect 2434 9998 2446 10001
rect 3154 9998 3166 10001
rect 3218 9998 3230 10050
rect 10446 9986 10498 9998
rect 12574 10050 12626 10062
rect 12574 9986 12626 9998
rect 17614 10050 17666 10062
rect 17614 9986 17666 9998
rect 19518 10050 19570 10062
rect 19518 9986 19570 9998
rect 21646 10050 21698 10062
rect 21646 9986 21698 9998
rect 30270 10050 30322 10062
rect 30270 9986 30322 9998
rect 36654 10050 36706 10062
rect 36654 9986 36706 9998
rect 37662 10050 37714 10062
rect 37662 9986 37714 9998
rect 2382 9938 2434 9950
rect 2382 9874 2434 9886
rect 2830 9938 2882 9950
rect 2830 9874 2882 9886
rect 4510 9938 4562 9950
rect 4510 9874 4562 9886
rect 5070 9938 5122 9950
rect 10334 9938 10386 9950
rect 19406 9938 19458 9950
rect 20862 9938 20914 9950
rect 24670 9938 24722 9950
rect 6626 9886 6638 9938
rect 6690 9886 6702 9938
rect 13682 9886 13694 9938
rect 13746 9886 13758 9938
rect 20626 9886 20638 9938
rect 20690 9886 20702 9938
rect 22530 9886 22542 9938
rect 22594 9886 22606 9938
rect 5070 9874 5122 9886
rect 10334 9874 10386 9886
rect 19406 9874 19458 9886
rect 20862 9874 20914 9886
rect 24670 9874 24722 9886
rect 25454 9938 25506 9950
rect 25454 9874 25506 9886
rect 27694 9938 27746 9950
rect 27694 9874 27746 9886
rect 30046 9938 30098 9950
rect 30046 9874 30098 9886
rect 30606 9938 30658 9950
rect 36766 9938 36818 9950
rect 39678 9938 39730 9950
rect 33170 9886 33182 9938
rect 33234 9886 33246 9938
rect 35298 9886 35310 9938
rect 35362 9886 35374 9938
rect 38770 9886 38782 9938
rect 38834 9886 38846 9938
rect 30606 9874 30658 9886
rect 36766 9874 36818 9886
rect 39678 9874 39730 9886
rect 11118 9826 11170 9838
rect 9426 9774 9438 9826
rect 9490 9774 9502 9826
rect 11118 9762 11170 9774
rect 11566 9826 11618 9838
rect 11566 9762 11618 9774
rect 11790 9826 11842 9838
rect 17278 9826 17330 9838
rect 16482 9774 16494 9826
rect 16546 9774 16558 9826
rect 11790 9762 11842 9774
rect 17278 9762 17330 9774
rect 17502 9826 17554 9838
rect 17502 9762 17554 9774
rect 18286 9826 18338 9838
rect 18286 9762 18338 9774
rect 19070 9826 19122 9838
rect 19070 9762 19122 9774
rect 19182 9826 19234 9838
rect 19182 9762 19234 9774
rect 21758 9826 21810 9838
rect 26014 9826 26066 9838
rect 22306 9774 22318 9826
rect 22370 9774 22382 9826
rect 22642 9774 22654 9826
rect 22706 9774 22718 9826
rect 23762 9774 23774 9826
rect 23826 9774 23838 9826
rect 21758 9762 21810 9774
rect 26014 9762 26066 9774
rect 26686 9826 26738 9838
rect 26686 9762 26738 9774
rect 27358 9826 27410 9838
rect 38558 9826 38610 9838
rect 28802 9774 28814 9826
rect 28866 9774 28878 9826
rect 31378 9774 31390 9826
rect 31442 9774 31454 9826
rect 31602 9774 31614 9826
rect 31666 9774 31678 9826
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 37538 9774 37550 9826
rect 37602 9774 37614 9826
rect 37762 9774 37774 9826
rect 37826 9774 37838 9826
rect 27358 9762 27410 9774
rect 38558 9762 38610 9774
rect 39790 9826 39842 9838
rect 39790 9762 39842 9774
rect 40910 9826 40962 9838
rect 40910 9762 40962 9774
rect 6078 9714 6130 9726
rect 12798 9714 12850 9726
rect 17166 9714 17218 9726
rect 8754 9662 8766 9714
rect 8818 9662 8830 9714
rect 15810 9662 15822 9714
rect 15874 9662 15886 9714
rect 6078 9650 6130 9662
rect 12798 9650 12850 9662
rect 17166 9650 17218 9662
rect 21982 9714 22034 9726
rect 21982 9650 22034 9662
rect 23998 9714 24050 9726
rect 23998 9650 24050 9662
rect 24558 9714 24610 9726
rect 24558 9650 24610 9662
rect 25006 9714 25058 9726
rect 25006 9650 25058 9662
rect 27470 9714 27522 9726
rect 27470 9650 27522 9662
rect 27806 9714 27858 9726
rect 27806 9650 27858 9662
rect 31166 9714 31218 9726
rect 31166 9650 31218 9662
rect 35982 9714 36034 9726
rect 35982 9650 36034 9662
rect 36094 9714 36146 9726
rect 36094 9650 36146 9662
rect 37998 9714 38050 9726
rect 37998 9650 38050 9662
rect 39566 9714 39618 9726
rect 39566 9650 39618 9662
rect 40126 9714 40178 9726
rect 40126 9650 40178 9662
rect 40574 9714 40626 9726
rect 40574 9650 40626 9662
rect 40798 9714 40850 9726
rect 40798 9650 40850 9662
rect 41694 9714 41746 9726
rect 41694 9650 41746 9662
rect 1934 9602 1986 9614
rect 1934 9538 1986 9550
rect 3166 9602 3218 9614
rect 3166 9538 3218 9550
rect 3614 9602 3666 9614
rect 3614 9538 3666 9550
rect 4174 9602 4226 9614
rect 4174 9538 4226 9550
rect 5630 9602 5682 9614
rect 5630 9538 5682 9550
rect 10222 9602 10274 9614
rect 10222 9538 10274 9550
rect 11454 9602 11506 9614
rect 11454 9538 11506 9550
rect 12686 9602 12738 9614
rect 12686 9538 12738 9550
rect 18398 9602 18450 9614
rect 18398 9538 18450 9550
rect 18622 9602 18674 9614
rect 18622 9538 18674 9550
rect 23438 9602 23490 9614
rect 23438 9538 23490 9550
rect 23550 9602 23602 9614
rect 23550 9538 23602 9550
rect 24782 9602 24834 9614
rect 24782 9538 24834 9550
rect 26462 9602 26514 9614
rect 26462 9538 26514 9550
rect 26574 9602 26626 9614
rect 26574 9538 26626 9550
rect 28254 9602 28306 9614
rect 28254 9538 28306 9550
rect 28366 9602 28418 9614
rect 28366 9538 28418 9550
rect 28590 9602 28642 9614
rect 28590 9538 28642 9550
rect 29486 9602 29538 9614
rect 29486 9538 29538 9550
rect 31054 9602 31106 9614
rect 31054 9538 31106 9550
rect 35758 9602 35810 9614
rect 35758 9538 35810 9550
rect 38782 9602 38834 9614
rect 38782 9538 38834 9550
rect 41358 9602 41410 9614
rect 41358 9538 41410 9550
rect 41582 9602 41634 9614
rect 41582 9538 41634 9550
rect 1344 9434 42560 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 42560 9434
rect 1344 9348 42560 9382
rect 3838 9266 3890 9278
rect 3838 9202 3890 9214
rect 7982 9266 8034 9278
rect 7982 9202 8034 9214
rect 9886 9266 9938 9278
rect 9886 9202 9938 9214
rect 10894 9266 10946 9278
rect 10894 9202 10946 9214
rect 17726 9266 17778 9278
rect 17726 9202 17778 9214
rect 18286 9266 18338 9278
rect 18286 9202 18338 9214
rect 24558 9266 24610 9278
rect 24558 9202 24610 9214
rect 25566 9266 25618 9278
rect 25566 9202 25618 9214
rect 25678 9266 25730 9278
rect 25678 9202 25730 9214
rect 25902 9266 25954 9278
rect 25902 9202 25954 9214
rect 26910 9266 26962 9278
rect 26910 9202 26962 9214
rect 27134 9266 27186 9278
rect 27134 9202 27186 9214
rect 27246 9266 27298 9278
rect 27246 9202 27298 9214
rect 29710 9266 29762 9278
rect 29710 9202 29762 9214
rect 31054 9266 31106 9278
rect 31054 9202 31106 9214
rect 31278 9266 31330 9278
rect 31278 9202 31330 9214
rect 31838 9266 31890 9278
rect 31838 9202 31890 9214
rect 32062 9266 32114 9278
rect 32062 9202 32114 9214
rect 32734 9266 32786 9278
rect 32734 9202 32786 9214
rect 33854 9266 33906 9278
rect 33854 9202 33906 9214
rect 34638 9266 34690 9278
rect 34638 9202 34690 9214
rect 37326 9266 37378 9278
rect 37326 9202 37378 9214
rect 38110 9266 38162 9278
rect 38110 9202 38162 9214
rect 38894 9266 38946 9278
rect 38894 9202 38946 9214
rect 39454 9266 39506 9278
rect 39454 9202 39506 9214
rect 40462 9266 40514 9278
rect 40462 9202 40514 9214
rect 5406 9154 5458 9166
rect 5406 9090 5458 9102
rect 5966 9154 6018 9166
rect 5966 9090 6018 9102
rect 6078 9154 6130 9166
rect 6078 9090 6130 9102
rect 6862 9154 6914 9166
rect 6862 9090 6914 9102
rect 7086 9154 7138 9166
rect 7086 9090 7138 9102
rect 7534 9154 7586 9166
rect 7534 9090 7586 9102
rect 8878 9154 8930 9166
rect 8878 9090 8930 9102
rect 10110 9154 10162 9166
rect 18510 9154 18562 9166
rect 11890 9102 11902 9154
rect 11954 9102 11966 9154
rect 10110 9090 10162 9102
rect 18510 9090 18562 9102
rect 26126 9154 26178 9166
rect 26126 9090 26178 9102
rect 26686 9154 26738 9166
rect 26686 9090 26738 9102
rect 27806 9154 27858 9166
rect 27806 9090 27858 9102
rect 28590 9154 28642 9166
rect 28590 9090 28642 9102
rect 29038 9154 29090 9166
rect 29038 9090 29090 9102
rect 29598 9154 29650 9166
rect 29598 9090 29650 9102
rect 30830 9154 30882 9166
rect 39678 9154 39730 9166
rect 36642 9102 36654 9154
rect 36706 9102 36718 9154
rect 30830 9090 30882 9102
rect 39678 9090 39730 9102
rect 39790 9154 39842 9166
rect 39790 9090 39842 9102
rect 40574 9154 40626 9166
rect 40574 9090 40626 9102
rect 41694 9154 41746 9166
rect 41694 9090 41746 9102
rect 41806 9154 41858 9166
rect 41806 9090 41858 9102
rect 6302 9042 6354 9054
rect 6302 8978 6354 8990
rect 6750 9042 6802 9054
rect 6750 8978 6802 8990
rect 7758 9042 7810 9054
rect 7758 8978 7810 8990
rect 8206 9042 8258 9054
rect 22990 9042 23042 9054
rect 16706 8990 16718 9042
rect 16770 8990 16782 9042
rect 22418 8990 22430 9042
rect 22482 8990 22494 9042
rect 8206 8978 8258 8990
rect 22990 8978 23042 8990
rect 23438 9042 23490 9054
rect 23438 8978 23490 8990
rect 23550 9042 23602 9054
rect 23550 8978 23602 8990
rect 23662 9042 23714 9054
rect 23662 8978 23714 8990
rect 24110 9042 24162 9054
rect 24110 8978 24162 8990
rect 24782 9042 24834 9054
rect 24782 8978 24834 8990
rect 27918 9042 27970 9054
rect 27918 8978 27970 8990
rect 28478 9042 28530 9054
rect 28478 8978 28530 8990
rect 28814 9042 28866 9054
rect 31390 9042 31442 9054
rect 34750 9042 34802 9054
rect 37438 9042 37490 9054
rect 29922 8990 29934 9042
rect 29986 8990 29998 9042
rect 32274 8990 32286 9042
rect 32338 8990 32350 9042
rect 35410 8990 35422 9042
rect 35474 8990 35486 9042
rect 28814 8978 28866 8990
rect 31390 8978 31442 8990
rect 34750 8978 34802 8990
rect 37438 8978 37490 8990
rect 37998 9042 38050 9054
rect 37998 8978 38050 8990
rect 39006 9042 39058 9054
rect 39006 8978 39058 8990
rect 41470 9042 41522 9054
rect 41470 8978 41522 8990
rect 2158 8930 2210 8942
rect 2158 8866 2210 8878
rect 2494 8930 2546 8942
rect 2494 8866 2546 8878
rect 3054 8930 3106 8942
rect 3054 8866 3106 8878
rect 3390 8930 3442 8942
rect 3390 8866 3442 8878
rect 4286 8930 4338 8942
rect 4286 8866 4338 8878
rect 4734 8930 4786 8942
rect 19182 8930 19234 8942
rect 24670 8930 24722 8942
rect 34862 8930 34914 8942
rect 36318 8930 36370 8942
rect 8978 8878 8990 8930
rect 9042 8878 9054 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 19618 8878 19630 8930
rect 19682 8878 19694 8930
rect 21746 8878 21758 8930
rect 21810 8878 21822 8930
rect 33954 8878 33966 8930
rect 34018 8878 34030 8930
rect 35522 8878 35534 8930
rect 35586 8878 35598 8930
rect 4734 8866 4786 8878
rect 19182 8866 19234 8878
rect 24670 8866 24722 8878
rect 34862 8866 34914 8878
rect 36318 8866 36370 8878
rect 5294 8818 5346 8830
rect 3378 8766 3390 8818
rect 3442 8815 3454 8818
rect 4498 8815 4510 8818
rect 3442 8769 4510 8815
rect 3442 8766 3454 8769
rect 4498 8766 4510 8769
rect 4562 8766 4574 8818
rect 5294 8754 5346 8766
rect 8654 8818 8706 8830
rect 8654 8754 8706 8766
rect 9774 8818 9826 8830
rect 9774 8754 9826 8766
rect 10670 8818 10722 8830
rect 10670 8754 10722 8766
rect 11006 8818 11058 8830
rect 11006 8754 11058 8766
rect 27806 8818 27858 8830
rect 27806 8754 27858 8766
rect 31726 8818 31778 8830
rect 31726 8754 31778 8766
rect 33630 8818 33682 8830
rect 33630 8754 33682 8766
rect 35758 8818 35810 8830
rect 35758 8754 35810 8766
rect 37326 8818 37378 8830
rect 37326 8754 37378 8766
rect 38110 8818 38162 8830
rect 38110 8754 38162 8766
rect 38894 8818 38946 8830
rect 38894 8754 38946 8766
rect 40462 8818 40514 8830
rect 40462 8754 40514 8766
rect 1344 8650 42560 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 42560 8650
rect 1344 8564 42560 8598
rect 6526 8482 6578 8494
rect 3378 8430 3390 8482
rect 3442 8479 3454 8482
rect 4050 8479 4062 8482
rect 3442 8433 4062 8479
rect 3442 8430 3454 8433
rect 4050 8430 4062 8433
rect 4114 8430 4126 8482
rect 6526 8418 6578 8430
rect 19630 8482 19682 8494
rect 19630 8418 19682 8430
rect 38446 8482 38498 8494
rect 38446 8418 38498 8430
rect 41694 8482 41746 8494
rect 41694 8418 41746 8430
rect 3390 8370 3442 8382
rect 3390 8306 3442 8318
rect 3838 8370 3890 8382
rect 3838 8306 3890 8318
rect 8542 8370 8594 8382
rect 14142 8370 14194 8382
rect 9986 8318 9998 8370
rect 10050 8318 10062 8370
rect 12114 8318 12126 8370
rect 12178 8318 12190 8370
rect 8542 8306 8594 8318
rect 14142 8306 14194 8318
rect 15150 8370 15202 8382
rect 20526 8370 20578 8382
rect 22094 8370 22146 8382
rect 28702 8370 28754 8382
rect 16818 8318 16830 8370
rect 16882 8318 16894 8370
rect 18946 8318 18958 8370
rect 19010 8318 19022 8370
rect 20738 8318 20750 8370
rect 20802 8318 20814 8370
rect 25218 8318 25230 8370
rect 25282 8318 25294 8370
rect 15150 8306 15202 8318
rect 20526 8306 20578 8318
rect 22094 8306 22146 8318
rect 28702 8306 28754 8318
rect 29598 8370 29650 8382
rect 30494 8370 30546 8382
rect 29810 8318 29822 8370
rect 29874 8318 29886 8370
rect 29598 8306 29650 8318
rect 30494 8306 30546 8318
rect 31390 8370 31442 8382
rect 36430 8370 36482 8382
rect 31714 8318 31726 8370
rect 31778 8318 31790 8370
rect 33394 8318 33406 8370
rect 33458 8318 33470 8370
rect 35522 8318 35534 8370
rect 35586 8318 35598 8370
rect 40674 8318 40686 8370
rect 40738 8318 40750 8370
rect 31390 8306 31442 8318
rect 36430 8306 36482 8318
rect 1934 8258 1986 8270
rect 1934 8194 1986 8206
rect 4174 8258 4226 8270
rect 4174 8194 4226 8206
rect 4734 8258 4786 8270
rect 4734 8194 4786 8206
rect 5966 8258 6018 8270
rect 5966 8194 6018 8206
rect 7758 8258 7810 8270
rect 14590 8258 14642 8270
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 8754 8206 8766 8258
rect 8818 8255 8830 8258
rect 8978 8255 8990 8258
rect 8818 8209 8990 8255
rect 8818 8206 8830 8209
rect 8978 8206 8990 8209
rect 9042 8206 9054 8258
rect 9426 8206 9438 8258
rect 9490 8206 9502 8258
rect 12786 8206 12798 8258
rect 12850 8206 12862 8258
rect 7758 8194 7810 8206
rect 14590 8194 14642 8206
rect 15038 8258 15090 8270
rect 15038 8194 15090 8206
rect 15262 8258 15314 8270
rect 22318 8258 22370 8270
rect 36542 8258 36594 8270
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 19954 8206 19966 8258
rect 20018 8206 20030 8258
rect 23874 8206 23886 8258
rect 23938 8206 23950 8258
rect 32610 8206 32622 8258
rect 32674 8206 32686 8258
rect 36082 8206 36094 8258
rect 36146 8206 36158 8258
rect 15262 8194 15314 8206
rect 22318 8194 22370 8206
rect 36542 8194 36594 8206
rect 37438 8258 37490 8270
rect 37438 8194 37490 8206
rect 38782 8258 38834 8270
rect 38782 8194 38834 8206
rect 39454 8258 39506 8270
rect 39454 8194 39506 8206
rect 39790 8258 39842 8270
rect 39790 8194 39842 8206
rect 5630 8146 5682 8158
rect 5630 8082 5682 8094
rect 6862 8146 6914 8158
rect 6862 8082 6914 8094
rect 7422 8146 7474 8158
rect 7422 8082 7474 8094
rect 9102 8146 9154 8158
rect 9102 8082 9154 8094
rect 13918 8146 13970 8158
rect 13918 8082 13970 8094
rect 21758 8146 21810 8158
rect 21758 8082 21810 8094
rect 22206 8146 22258 8158
rect 22206 8082 22258 8094
rect 36766 8146 36818 8158
rect 36766 8082 36818 8094
rect 37662 8146 37714 8158
rect 37662 8082 37714 8094
rect 37774 8146 37826 8158
rect 37774 8082 37826 8094
rect 39006 8146 39058 8158
rect 39006 8082 39058 8094
rect 40126 8146 40178 8158
rect 40126 8082 40178 8094
rect 41022 8146 41074 8158
rect 41022 8082 41074 8094
rect 41694 8146 41746 8158
rect 41694 8082 41746 8094
rect 41806 8146 41858 8158
rect 41806 8082 41858 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 2830 8034 2882 8046
rect 2830 7970 2882 7982
rect 4846 8034 4898 8046
rect 4846 7970 4898 7982
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 5854 8034 5906 8046
rect 5854 7970 5906 7982
rect 6638 8034 6690 8046
rect 6638 7970 6690 7982
rect 7534 8034 7586 8046
rect 7534 7970 7586 7982
rect 8430 8034 8482 8046
rect 8430 7970 8482 7982
rect 9214 8034 9266 8046
rect 9214 7970 9266 7982
rect 14030 8034 14082 8046
rect 14030 7970 14082 7982
rect 19742 8034 19794 8046
rect 19742 7970 19794 7982
rect 21982 8034 22034 8046
rect 21982 7970 22034 7982
rect 29822 8034 29874 8046
rect 29822 7970 29874 7982
rect 30606 8034 30658 8046
rect 30606 7970 30658 7982
rect 31614 8034 31666 8046
rect 31614 7970 31666 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 39790 8034 39842 8046
rect 39790 7970 39842 7982
rect 1344 7866 42560 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 42560 7866
rect 1344 7780 42560 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 2270 7698 2322 7710
rect 2270 7634 2322 7646
rect 2718 7698 2770 7710
rect 2718 7634 2770 7646
rect 3054 7698 3106 7710
rect 3054 7634 3106 7646
rect 6750 7698 6802 7710
rect 6750 7634 6802 7646
rect 7870 7698 7922 7710
rect 7870 7634 7922 7646
rect 8878 7698 8930 7710
rect 8878 7634 8930 7646
rect 10334 7698 10386 7710
rect 10334 7634 10386 7646
rect 10558 7698 10610 7710
rect 10558 7634 10610 7646
rect 21310 7698 21362 7710
rect 21310 7634 21362 7646
rect 23102 7698 23154 7710
rect 23102 7634 23154 7646
rect 25566 7698 25618 7710
rect 29710 7698 29762 7710
rect 26786 7646 26798 7698
rect 26850 7646 26862 7698
rect 25566 7634 25618 7646
rect 29710 7634 29762 7646
rect 30606 7698 30658 7710
rect 30606 7634 30658 7646
rect 31726 7698 31778 7710
rect 31726 7634 31778 7646
rect 33742 7698 33794 7710
rect 33742 7634 33794 7646
rect 35646 7698 35698 7710
rect 37886 7698 37938 7710
rect 36642 7646 36654 7698
rect 36706 7646 36718 7698
rect 35646 7634 35698 7646
rect 37886 7634 37938 7646
rect 37998 7698 38050 7710
rect 37998 7634 38050 7646
rect 38222 7698 38274 7710
rect 38222 7634 38274 7646
rect 39118 7698 39170 7710
rect 39118 7634 39170 7646
rect 40014 7698 40066 7710
rect 40014 7634 40066 7646
rect 41694 7698 41746 7710
rect 41694 7634 41746 7646
rect 3726 7586 3778 7598
rect 3726 7522 3778 7534
rect 4286 7586 4338 7598
rect 4286 7522 4338 7534
rect 4958 7586 5010 7598
rect 4958 7522 5010 7534
rect 5070 7586 5122 7598
rect 5070 7522 5122 7534
rect 5854 7586 5906 7598
rect 5854 7522 5906 7534
rect 6974 7586 7026 7598
rect 6974 7522 7026 7534
rect 10110 7586 10162 7598
rect 10110 7522 10162 7534
rect 21198 7586 21250 7598
rect 21198 7522 21250 7534
rect 21422 7586 21474 7598
rect 22430 7586 22482 7598
rect 22082 7534 22094 7586
rect 22146 7534 22158 7586
rect 21422 7522 21474 7534
rect 22430 7522 22482 7534
rect 23886 7586 23938 7598
rect 23886 7522 23938 7534
rect 26238 7586 26290 7598
rect 26238 7522 26290 7534
rect 27918 7586 27970 7598
rect 35534 7586 35586 7598
rect 32498 7534 32510 7586
rect 32562 7534 32574 7586
rect 27918 7522 27970 7534
rect 35534 7522 35586 7534
rect 36094 7586 36146 7598
rect 36094 7522 36146 7534
rect 39342 7586 39394 7598
rect 39342 7522 39394 7534
rect 39902 7586 39954 7598
rect 39902 7522 39954 7534
rect 41806 7586 41858 7598
rect 41806 7522 41858 7534
rect 4398 7474 4450 7486
rect 4398 7410 4450 7422
rect 5294 7474 5346 7486
rect 5294 7410 5346 7422
rect 5742 7474 5794 7486
rect 5742 7410 5794 7422
rect 6638 7474 6690 7486
rect 6638 7410 6690 7422
rect 7086 7474 7138 7486
rect 7086 7410 7138 7422
rect 8542 7474 8594 7486
rect 8542 7410 8594 7422
rect 8766 7474 8818 7486
rect 10670 7474 10722 7486
rect 22990 7474 23042 7486
rect 26462 7474 26514 7486
rect 28478 7474 28530 7486
rect 8978 7422 8990 7474
rect 9042 7422 9054 7474
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 17826 7422 17838 7474
rect 17890 7422 17902 7474
rect 23650 7422 23662 7474
rect 23714 7422 23726 7474
rect 27458 7422 27470 7474
rect 27522 7422 27534 7474
rect 8766 7410 8818 7422
rect 10670 7410 10722 7422
rect 22990 7410 23042 7422
rect 26462 7410 26514 7422
rect 28478 7410 28530 7422
rect 28814 7474 28866 7486
rect 28814 7410 28866 7422
rect 29038 7474 29090 7486
rect 29038 7410 29090 7422
rect 30494 7474 30546 7486
rect 31838 7474 31890 7486
rect 30818 7422 30830 7474
rect 30882 7422 30894 7474
rect 30494 7410 30546 7422
rect 31838 7410 31890 7422
rect 32846 7474 32898 7486
rect 32846 7410 32898 7422
rect 34526 7474 34578 7486
rect 38558 7474 38610 7486
rect 34850 7422 34862 7474
rect 34914 7422 34926 7474
rect 36754 7422 36766 7474
rect 36818 7422 36830 7474
rect 36978 7422 36990 7474
rect 37042 7422 37054 7474
rect 40226 7422 40238 7474
rect 40290 7422 40302 7474
rect 34526 7410 34578 7422
rect 38558 7410 38610 7422
rect 3614 7362 3666 7374
rect 3614 7298 3666 7310
rect 6862 7362 6914 7374
rect 6862 7298 6914 7310
rect 7758 7362 7810 7374
rect 23214 7362 23266 7374
rect 11778 7310 11790 7362
rect 11842 7310 11854 7362
rect 18498 7310 18510 7362
rect 18562 7310 18574 7362
rect 20626 7310 20638 7362
rect 20690 7310 20702 7362
rect 7758 7298 7810 7310
rect 23214 7298 23266 7310
rect 24446 7362 24498 7374
rect 28590 7362 28642 7374
rect 31278 7362 31330 7374
rect 24658 7310 24670 7362
rect 24722 7310 24734 7362
rect 29586 7310 29598 7362
rect 29650 7310 29662 7362
rect 24446 7298 24498 7310
rect 28590 7298 28642 7310
rect 31278 7298 31330 7310
rect 32062 7362 32114 7374
rect 35310 7362 35362 7374
rect 33618 7310 33630 7362
rect 33682 7310 33694 7362
rect 32062 7298 32114 7310
rect 35310 7298 35362 7310
rect 36318 7362 36370 7374
rect 36318 7298 36370 7310
rect 37438 7362 37490 7374
rect 37438 7298 37490 7310
rect 39230 7362 39282 7374
rect 39230 7298 39282 7310
rect 40686 7362 40738 7374
rect 40686 7298 40738 7310
rect 5854 7250 5906 7262
rect 5854 7186 5906 7198
rect 10222 7250 10274 7262
rect 10222 7186 10274 7198
rect 23438 7250 23490 7262
rect 23438 7186 23490 7198
rect 29934 7250 29986 7262
rect 29934 7186 29986 7198
rect 32286 7250 32338 7262
rect 32286 7186 32338 7198
rect 33966 7250 34018 7262
rect 33966 7186 34018 7198
rect 35086 7250 35138 7262
rect 35086 7186 35138 7198
rect 36542 7250 36594 7262
rect 36542 7186 36594 7198
rect 41694 7250 41746 7262
rect 41694 7186 41746 7198
rect 1344 7082 42560 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 42560 7082
rect 1344 6996 42560 7030
rect 17278 6914 17330 6926
rect 17278 6850 17330 6862
rect 24110 6914 24162 6926
rect 24110 6850 24162 6862
rect 1934 6802 1986 6814
rect 6514 6750 6526 6802
rect 6578 6750 6590 6802
rect 9986 6750 9998 6802
rect 10050 6750 10062 6802
rect 16818 6750 16830 6802
rect 16882 6750 16894 6802
rect 35074 6750 35086 6802
rect 35138 6750 35150 6802
rect 38994 6750 39006 6802
rect 39058 6750 39070 6802
rect 1934 6738 1986 6750
rect 2382 6690 2434 6702
rect 2382 6626 2434 6638
rect 3278 6690 3330 6702
rect 18622 6690 18674 6702
rect 19406 6690 19458 6702
rect 8642 6638 8654 6690
rect 8706 6638 8718 6690
rect 9426 6638 9438 6690
rect 9490 6638 9502 6690
rect 12786 6638 12798 6690
rect 12850 6638 12862 6690
rect 13906 6638 13918 6690
rect 13970 6638 13982 6690
rect 18946 6638 18958 6690
rect 19010 6638 19022 6690
rect 3278 6626 3330 6638
rect 18622 6626 18674 6638
rect 19406 6626 19458 6638
rect 19854 6690 19906 6702
rect 19854 6626 19906 6638
rect 20638 6690 20690 6702
rect 20638 6626 20690 6638
rect 20974 6690 21026 6702
rect 23214 6690 23266 6702
rect 25454 6690 25506 6702
rect 22754 6638 22766 6690
rect 22818 6638 22830 6690
rect 23426 6638 23438 6690
rect 23490 6638 23502 6690
rect 20974 6626 21026 6638
rect 23214 6626 23266 6638
rect 25454 6626 25506 6638
rect 25678 6690 25730 6702
rect 26350 6690 26402 6702
rect 25890 6638 25902 6690
rect 25954 6638 25966 6690
rect 25678 6626 25730 6638
rect 26350 6626 26402 6638
rect 27022 6690 27074 6702
rect 27022 6626 27074 6638
rect 28142 6690 28194 6702
rect 28142 6626 28194 6638
rect 28702 6690 28754 6702
rect 28702 6626 28754 6638
rect 28814 6690 28866 6702
rect 28814 6626 28866 6638
rect 30158 6690 30210 6702
rect 31390 6690 31442 6702
rect 38446 6690 38498 6702
rect 30370 6638 30382 6690
rect 30434 6638 30446 6690
rect 31602 6638 31614 6690
rect 31666 6638 31678 6690
rect 32274 6638 32286 6690
rect 32338 6638 32350 6690
rect 36642 6638 36654 6690
rect 36706 6638 36718 6690
rect 30158 6626 30210 6638
rect 31390 6626 31442 6638
rect 38446 6626 38498 6638
rect 40910 6690 40962 6702
rect 40910 6626 40962 6638
rect 41582 6690 41634 6702
rect 41582 6626 41634 6638
rect 41918 6690 41970 6702
rect 41918 6626 41970 6638
rect 4174 6578 4226 6590
rect 4174 6514 4226 6526
rect 4846 6578 4898 6590
rect 4846 6514 4898 6526
rect 5966 6578 6018 6590
rect 17390 6578 17442 6590
rect 12114 6526 12126 6578
rect 12178 6526 12190 6578
rect 14690 6526 14702 6578
rect 14754 6526 14766 6578
rect 5966 6514 6018 6526
rect 17390 6514 17442 6526
rect 17838 6578 17890 6590
rect 17838 6514 17890 6526
rect 20078 6578 20130 6590
rect 20078 6514 20130 6526
rect 21646 6578 21698 6590
rect 21646 6514 21698 6526
rect 22206 6578 22258 6590
rect 22206 6514 22258 6526
rect 23998 6578 24050 6590
rect 23998 6514 24050 6526
rect 24670 6578 24722 6590
rect 24670 6514 24722 6526
rect 25230 6578 25282 6590
rect 25230 6514 25282 6526
rect 26798 6578 26850 6590
rect 26798 6514 26850 6526
rect 27694 6578 27746 6590
rect 27694 6514 27746 6526
rect 29710 6578 29762 6590
rect 29710 6514 29762 6526
rect 30942 6578 30994 6590
rect 30942 6514 30994 6526
rect 31278 6578 31330 6590
rect 35982 6578 36034 6590
rect 32946 6526 32958 6578
rect 33010 6526 33022 6578
rect 31278 6514 31330 6526
rect 35982 6514 36034 6526
rect 37886 6578 37938 6590
rect 41022 6578 41074 6590
rect 39890 6526 39902 6578
rect 39954 6526 39966 6578
rect 37886 6514 37938 6526
rect 41022 6514 41074 6526
rect 41806 6578 41858 6590
rect 41806 6514 41858 6526
rect 2718 6466 2770 6478
rect 2718 6402 2770 6414
rect 3726 6466 3778 6478
rect 3726 6402 3778 6414
rect 4286 6466 4338 6478
rect 4286 6402 4338 6414
rect 4958 6466 5010 6478
rect 4958 6402 5010 6414
rect 5630 6466 5682 6478
rect 5630 6402 5682 6414
rect 5854 6466 5906 6478
rect 5854 6402 5906 6414
rect 17614 6466 17666 6478
rect 17614 6402 17666 6414
rect 18398 6466 18450 6478
rect 18398 6402 18450 6414
rect 18510 6466 18562 6478
rect 18510 6402 18562 6414
rect 19630 6466 19682 6478
rect 19630 6402 19682 6414
rect 20750 6466 20802 6478
rect 20750 6402 20802 6414
rect 22990 6466 23042 6478
rect 22990 6402 23042 6414
rect 23102 6466 23154 6478
rect 23102 6402 23154 6414
rect 24222 6466 24274 6478
rect 24222 6402 24274 6414
rect 24446 6466 24498 6478
rect 24446 6402 24498 6414
rect 25566 6466 25618 6478
rect 25566 6402 25618 6414
rect 26686 6466 26738 6478
rect 26686 6402 26738 6414
rect 27918 6466 27970 6478
rect 27918 6402 27970 6414
rect 28030 6466 28082 6478
rect 28030 6402 28082 6414
rect 29934 6466 29986 6478
rect 29934 6402 29986 6414
rect 30046 6466 30098 6478
rect 30046 6402 30098 6414
rect 31166 6466 31218 6478
rect 31166 6402 31218 6414
rect 36206 6466 36258 6478
rect 36206 6402 36258 6414
rect 36318 6466 36370 6478
rect 36318 6402 36370 6414
rect 36430 6466 36482 6478
rect 36430 6402 36482 6414
rect 37774 6466 37826 6478
rect 37774 6402 37826 6414
rect 38110 6466 38162 6478
rect 38110 6402 38162 6414
rect 41246 6466 41298 6478
rect 41246 6402 41298 6414
rect 1344 6298 42560 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 42560 6298
rect 1344 6212 42560 6246
rect 2270 6130 2322 6142
rect 2270 6066 2322 6078
rect 2718 6130 2770 6142
rect 2718 6066 2770 6078
rect 3166 6130 3218 6142
rect 3166 6066 3218 6078
rect 4622 6130 4674 6142
rect 4622 6066 4674 6078
rect 6750 6130 6802 6142
rect 6750 6066 6802 6078
rect 9774 6130 9826 6142
rect 9774 6066 9826 6078
rect 10334 6130 10386 6142
rect 10334 6066 10386 6078
rect 10446 6130 10498 6142
rect 10446 6066 10498 6078
rect 11566 6130 11618 6142
rect 11566 6066 11618 6078
rect 14030 6130 14082 6142
rect 14030 6066 14082 6078
rect 14702 6130 14754 6142
rect 14702 6066 14754 6078
rect 16606 6130 16658 6142
rect 16606 6066 16658 6078
rect 16830 6130 16882 6142
rect 16830 6066 16882 6078
rect 19854 6130 19906 6142
rect 19854 6066 19906 6078
rect 23662 6130 23714 6142
rect 23662 6066 23714 6078
rect 25566 6130 25618 6142
rect 25566 6066 25618 6078
rect 26014 6130 26066 6142
rect 26014 6066 26066 6078
rect 27694 6130 27746 6142
rect 32734 6130 32786 6142
rect 30930 6078 30942 6130
rect 30994 6078 31006 6130
rect 27694 6066 27746 6078
rect 32734 6066 32786 6078
rect 37326 6130 37378 6142
rect 37326 6066 37378 6078
rect 37550 6130 37602 6142
rect 37550 6066 37602 6078
rect 38222 6130 38274 6142
rect 38222 6066 38274 6078
rect 40798 6130 40850 6142
rect 40798 6066 40850 6078
rect 41470 6130 41522 6142
rect 41470 6066 41522 6078
rect 41694 6130 41746 6142
rect 41694 6066 41746 6078
rect 5518 6018 5570 6030
rect 5518 5954 5570 5966
rect 5742 6018 5794 6030
rect 5742 5954 5794 5966
rect 6974 6018 7026 6030
rect 6974 5954 7026 5966
rect 8878 6018 8930 6030
rect 8878 5954 8930 5966
rect 11118 6018 11170 6030
rect 11118 5954 11170 5966
rect 11342 6018 11394 6030
rect 11342 5954 11394 5966
rect 11678 6018 11730 6030
rect 14814 6018 14866 6030
rect 12450 5966 12462 6018
rect 12514 5966 12526 6018
rect 13010 5966 13022 6018
rect 13074 5966 13086 6018
rect 11678 5954 11730 5966
rect 14814 5954 14866 5966
rect 15934 6018 15986 6030
rect 15934 5954 15986 5966
rect 16158 6018 16210 6030
rect 16158 5954 16210 5966
rect 16942 6018 16994 6030
rect 27022 6018 27074 6030
rect 37774 6018 37826 6030
rect 41806 6018 41858 6030
rect 17826 5966 17838 6018
rect 17890 5966 17902 6018
rect 22418 5966 22430 6018
rect 22482 5966 22494 6018
rect 29250 5966 29262 6018
rect 29314 5966 29326 6018
rect 40114 5966 40126 6018
rect 40178 5966 40190 6018
rect 16942 5954 16994 5966
rect 27022 5954 27074 5966
rect 37774 5954 37826 5966
rect 41806 5954 41858 5966
rect 4734 5906 4786 5918
rect 6526 5906 6578 5918
rect 6290 5854 6302 5906
rect 6354 5854 6366 5906
rect 4734 5842 4786 5854
rect 6526 5842 6578 5854
rect 8094 5906 8146 5918
rect 8094 5842 8146 5854
rect 12238 5906 12290 5918
rect 12238 5842 12290 5854
rect 14478 5906 14530 5918
rect 14478 5842 14530 5854
rect 15038 5906 15090 5918
rect 15038 5842 15090 5854
rect 15486 5906 15538 5918
rect 23774 5906 23826 5918
rect 17938 5854 17950 5906
rect 18002 5854 18014 5906
rect 18610 5854 18622 5906
rect 18674 5854 18686 5906
rect 19058 5854 19070 5906
rect 19122 5854 19134 5906
rect 23090 5854 23102 5906
rect 23154 5854 23166 5906
rect 15486 5842 15538 5854
rect 23774 5842 23826 5854
rect 23998 5906 24050 5918
rect 24782 5906 24834 5918
rect 24434 5854 24446 5906
rect 24498 5854 24510 5906
rect 23998 5842 24050 5854
rect 24782 5842 24834 5854
rect 26126 5906 26178 5918
rect 26126 5842 26178 5854
rect 26350 5906 26402 5918
rect 27582 5906 27634 5918
rect 26786 5854 26798 5906
rect 26850 5854 26862 5906
rect 26350 5842 26402 5854
rect 27582 5842 27634 5854
rect 30494 5906 30546 5918
rect 30494 5842 30546 5854
rect 30942 5906 30994 5918
rect 30942 5842 30994 5854
rect 31502 5906 31554 5918
rect 31502 5842 31554 5854
rect 32398 5906 32450 5918
rect 37214 5906 37266 5918
rect 36418 5854 36430 5906
rect 36482 5854 36494 5906
rect 32398 5842 32450 5854
rect 37214 5842 37266 5854
rect 1822 5794 1874 5806
rect 1822 5730 1874 5742
rect 3614 5794 3666 5806
rect 3614 5730 3666 5742
rect 4062 5794 4114 5806
rect 4062 5730 4114 5742
rect 6638 5794 6690 5806
rect 6638 5730 6690 5742
rect 8318 5794 8370 5806
rect 8318 5730 8370 5742
rect 12126 5794 12178 5806
rect 12126 5730 12178 5742
rect 15710 5794 15762 5806
rect 31054 5794 31106 5806
rect 20290 5742 20302 5794
rect 20354 5742 20366 5794
rect 28242 5742 28254 5794
rect 28306 5742 28318 5794
rect 15710 5730 15762 5742
rect 31054 5730 31106 5742
rect 31278 5794 31330 5806
rect 37438 5794 37490 5806
rect 33618 5742 33630 5794
rect 33682 5742 33694 5794
rect 35746 5742 35758 5794
rect 35810 5742 35822 5794
rect 38882 5742 38894 5794
rect 38946 5742 38958 5794
rect 31278 5730 31330 5742
rect 37438 5730 37490 5742
rect 4846 5682 4898 5694
rect 2146 5630 2158 5682
rect 2210 5679 2222 5682
rect 2930 5679 2942 5682
rect 2210 5633 2942 5679
rect 2210 5630 2222 5633
rect 2930 5630 2942 5633
rect 2994 5630 3006 5682
rect 4846 5618 4898 5630
rect 5406 5682 5458 5694
rect 8990 5682 9042 5694
rect 7746 5630 7758 5682
rect 7810 5630 7822 5682
rect 5406 5618 5458 5630
rect 8990 5618 9042 5630
rect 10558 5682 10610 5694
rect 24222 5682 24274 5694
rect 18946 5630 18958 5682
rect 19010 5630 19022 5682
rect 10558 5618 10610 5630
rect 24222 5618 24274 5630
rect 26574 5682 26626 5694
rect 26574 5618 26626 5630
rect 32174 5682 32226 5694
rect 32174 5618 32226 5630
rect 32622 5682 32674 5694
rect 32622 5618 32674 5630
rect 32734 5682 32786 5694
rect 32734 5618 32786 5630
rect 1344 5514 42560 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 42560 5514
rect 1344 5428 42560 5462
rect 3950 5346 4002 5358
rect 3950 5282 4002 5294
rect 6078 5346 6130 5358
rect 6078 5282 6130 5294
rect 23662 5346 23714 5358
rect 23662 5282 23714 5294
rect 24222 5346 24274 5358
rect 24222 5282 24274 5294
rect 25006 5346 25058 5358
rect 25006 5282 25058 5294
rect 28366 5346 28418 5358
rect 28366 5282 28418 5294
rect 35758 5346 35810 5358
rect 35758 5282 35810 5294
rect 35870 5346 35922 5358
rect 35870 5282 35922 5294
rect 41806 5346 41858 5358
rect 41806 5282 41858 5294
rect 2158 5234 2210 5246
rect 2158 5170 2210 5182
rect 2606 5234 2658 5246
rect 2606 5170 2658 5182
rect 3166 5234 3218 5246
rect 3166 5170 3218 5182
rect 6302 5234 6354 5246
rect 10334 5234 10386 5246
rect 6850 5182 6862 5234
rect 6914 5182 6926 5234
rect 8978 5182 8990 5234
rect 9042 5182 9054 5234
rect 6302 5170 6354 5182
rect 10334 5170 10386 5182
rect 12910 5234 12962 5246
rect 12910 5170 12962 5182
rect 13806 5234 13858 5246
rect 20862 5234 20914 5246
rect 28590 5234 28642 5246
rect 15026 5182 15038 5234
rect 15090 5182 15102 5234
rect 17154 5182 17166 5234
rect 17218 5182 17230 5234
rect 18386 5182 18398 5234
rect 18450 5182 18462 5234
rect 22306 5182 22318 5234
rect 22370 5182 22382 5234
rect 25554 5182 25566 5234
rect 25618 5182 25630 5234
rect 31042 5182 31054 5234
rect 31106 5182 31118 5234
rect 31602 5182 31614 5234
rect 31666 5182 31678 5234
rect 33730 5182 33742 5234
rect 33794 5182 33806 5234
rect 37650 5182 37662 5234
rect 37714 5182 37726 5234
rect 39666 5182 39678 5234
rect 39730 5182 39742 5234
rect 13806 5170 13858 5182
rect 20862 5170 20914 5182
rect 28590 5170 28642 5182
rect 4062 5122 4114 5134
rect 12574 5122 12626 5134
rect 19854 5122 19906 5134
rect 23886 5122 23938 5134
rect 5730 5070 5742 5122
rect 5794 5070 5806 5122
rect 9650 5070 9662 5122
rect 9714 5070 9726 5122
rect 14242 5070 14254 5122
rect 14306 5070 14318 5122
rect 17714 5070 17726 5122
rect 17778 5070 17790 5122
rect 21746 5070 21758 5122
rect 21810 5070 21822 5122
rect 4062 5058 4114 5070
rect 12574 5058 12626 5070
rect 19854 5058 19906 5070
rect 23886 5058 23938 5070
rect 24110 5122 24162 5134
rect 24110 5058 24162 5070
rect 27806 5122 27858 5134
rect 27806 5058 27858 5070
rect 28814 5122 28866 5134
rect 28814 5058 28866 5070
rect 36094 5122 36146 5134
rect 36094 5058 36146 5070
rect 36318 5122 36370 5134
rect 36318 5058 36370 5070
rect 41918 5122 41970 5134
rect 41918 5058 41970 5070
rect 4622 5010 4674 5022
rect 4622 4946 4674 4958
rect 10782 5010 10834 5022
rect 10782 4946 10834 4958
rect 11118 5010 11170 5022
rect 11118 4946 11170 4958
rect 11342 5010 11394 5022
rect 11342 4946 11394 4958
rect 11902 5010 11954 5022
rect 11902 4946 11954 4958
rect 12014 5010 12066 5022
rect 12014 4946 12066 4958
rect 19518 5010 19570 5022
rect 19518 4946 19570 4958
rect 19630 5010 19682 5022
rect 19630 4946 19682 4958
rect 20302 5010 20354 5022
rect 20302 4946 20354 4958
rect 24894 5010 24946 5022
rect 41806 5010 41858 5022
rect 26562 4958 26574 5010
rect 26626 4958 26638 5010
rect 28130 4958 28142 5010
rect 28194 4958 28206 5010
rect 29698 4958 29710 5010
rect 29762 4958 29774 5010
rect 32610 4958 32622 5010
rect 32674 4958 32686 5010
rect 34962 4958 34974 5010
rect 35026 4958 35038 5010
rect 38882 4958 38894 5010
rect 38946 4958 38958 5010
rect 40674 4958 40686 5010
rect 40738 4958 40750 5010
rect 24894 4946 24946 4958
rect 41806 4946 41858 4958
rect 3054 4898 3106 4910
rect 3054 4834 3106 4846
rect 3950 4898 4002 4910
rect 3950 4834 4002 4846
rect 4958 4898 5010 4910
rect 4958 4834 5010 4846
rect 10894 4898 10946 4910
rect 10894 4834 10946 4846
rect 12126 4898 12178 4910
rect 12126 4834 12178 4846
rect 23774 4898 23826 4910
rect 36206 4898 36258 4910
rect 28242 4846 28254 4898
rect 28306 4846 28318 4898
rect 23774 4834 23826 4846
rect 36206 4834 36258 4846
rect 1344 4730 42560 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 42560 4730
rect 1344 4644 42560 4678
rect 4734 4562 4786 4574
rect 16830 4562 16882 4574
rect 14242 4510 14254 4562
rect 14306 4510 14318 4562
rect 4734 4498 4786 4510
rect 16830 4498 16882 4510
rect 24782 4562 24834 4574
rect 24782 4498 24834 4510
rect 25790 4562 25842 4574
rect 25790 4498 25842 4510
rect 26014 4562 26066 4574
rect 26014 4498 26066 4510
rect 3614 4450 3666 4462
rect 3614 4386 3666 4398
rect 3950 4450 4002 4462
rect 3950 4386 4002 4398
rect 4510 4450 4562 4462
rect 16606 4450 16658 4462
rect 25678 4450 25730 4462
rect 10546 4398 10558 4450
rect 10610 4398 10622 4450
rect 19954 4398 19966 4450
rect 20018 4398 20030 4450
rect 23426 4398 23438 4450
rect 23490 4398 23502 4450
rect 30706 4398 30718 4450
rect 30770 4398 30782 4450
rect 35746 4398 35758 4450
rect 35810 4398 35822 4450
rect 38434 4398 38446 4450
rect 38498 4398 38510 4450
rect 40114 4398 40126 4450
rect 40178 4398 40190 4450
rect 41570 4398 41582 4450
rect 41634 4398 41646 4450
rect 4510 4386 4562 4398
rect 16606 4386 16658 4398
rect 25678 4386 25730 4398
rect 13694 4338 13746 4350
rect 2930 4286 2942 4338
rect 2994 4286 3006 4338
rect 5394 4286 5406 4338
rect 5458 4286 5470 4338
rect 7746 4286 7758 4338
rect 7810 4286 7822 4338
rect 9762 4286 9774 4338
rect 9826 4286 9838 4338
rect 13694 4274 13746 4286
rect 13918 4338 13970 4350
rect 24894 4338 24946 4350
rect 14914 4286 14926 4338
rect 14978 4286 14990 4338
rect 20738 4286 20750 4338
rect 20802 4286 20814 4338
rect 24098 4286 24110 4338
rect 24162 4286 24174 4338
rect 26450 4286 26462 4338
rect 26514 4286 26526 4338
rect 29922 4286 29934 4338
rect 29986 4286 29998 4338
rect 36418 4286 36430 4338
rect 36482 4286 36494 4338
rect 41794 4286 41806 4338
rect 41858 4286 41870 4338
rect 13918 4274 13970 4286
rect 24894 4274 24946 4286
rect 7310 4226 7362 4238
rect 13246 4226 13298 4238
rect 1922 4174 1934 4226
rect 1986 4174 1998 4226
rect 6066 4174 6078 4226
rect 6130 4174 6142 4226
rect 8418 4174 8430 4226
rect 8482 4174 8494 4226
rect 12674 4174 12686 4226
rect 12738 4174 12750 4226
rect 15474 4174 15486 4226
rect 15538 4174 15550 4226
rect 16930 4174 16942 4226
rect 16994 4174 17006 4226
rect 17826 4174 17838 4226
rect 17890 4174 17902 4226
rect 21298 4174 21310 4226
rect 21362 4174 21374 4226
rect 27234 4174 27246 4226
rect 27298 4174 27310 4226
rect 29362 4174 29374 4226
rect 29426 4174 29438 4226
rect 32834 4174 32846 4226
rect 32898 4174 32910 4226
rect 33618 4174 33630 4226
rect 33682 4174 33694 4226
rect 37090 4174 37102 4226
rect 37154 4174 37166 4226
rect 39106 4174 39118 4226
rect 39170 4174 39182 4226
rect 7310 4162 7362 4174
rect 13246 4162 13298 4174
rect 4846 4114 4898 4126
rect 4846 4050 4898 4062
rect 1344 3946 42560 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 42560 3946
rect 1344 3860 42560 3894
rect 21422 3778 21474 3790
rect 21422 3714 21474 3726
rect 31950 3778 32002 3790
rect 31950 3714 32002 3726
rect 35534 3778 35586 3790
rect 35534 3714 35586 3726
rect 35758 3778 35810 3790
rect 35758 3714 35810 3726
rect 21534 3666 21586 3678
rect 2482 3614 2494 3666
rect 2546 3614 2558 3666
rect 6514 3614 6526 3666
rect 6578 3614 6590 3666
rect 10546 3614 10558 3666
rect 10610 3614 10622 3666
rect 12226 3614 12238 3666
rect 12290 3614 12302 3666
rect 14242 3614 14254 3666
rect 14306 3614 14318 3666
rect 16146 3614 16158 3666
rect 16210 3614 16222 3666
rect 18610 3614 18622 3666
rect 18674 3614 18686 3666
rect 20178 3614 20190 3666
rect 20242 3614 20254 3666
rect 21534 3602 21586 3614
rect 24334 3666 24386 3678
rect 27694 3666 27746 3678
rect 25330 3614 25342 3666
rect 25394 3614 25406 3666
rect 24334 3602 24386 3614
rect 27694 3602 27746 3614
rect 28590 3666 28642 3678
rect 32174 3666 32226 3678
rect 35870 3666 35922 3678
rect 42030 3666 42082 3678
rect 29250 3614 29262 3666
rect 29314 3614 29326 3666
rect 33170 3614 33182 3666
rect 33234 3614 33246 3666
rect 37090 3614 37102 3666
rect 37154 3614 37166 3666
rect 28590 3602 28642 3614
rect 32174 3602 32226 3614
rect 35870 3602 35922 3614
rect 42030 3602 42082 3614
rect 27582 3554 27634 3566
rect 3042 3502 3054 3554
rect 3106 3502 3118 3554
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 5842 3502 5854 3554
rect 5906 3502 5918 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 9762 3502 9774 3554
rect 9826 3502 9838 3554
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 13570 3502 13582 3554
rect 13634 3502 13646 3554
rect 15586 3502 15598 3554
rect 15650 3502 15662 3554
rect 17602 3502 17614 3554
rect 17666 3502 17678 3554
rect 19394 3502 19406 3554
rect 19458 3502 19470 3554
rect 27346 3502 27358 3554
rect 27410 3502 27422 3554
rect 27582 3490 27634 3502
rect 27806 3554 27858 3566
rect 31390 3554 31442 3566
rect 28018 3502 28030 3554
rect 28082 3502 28094 3554
rect 27806 3490 27858 3502
rect 31390 3490 31442 3502
rect 31838 3554 31890 3566
rect 31838 3490 31890 3502
rect 32398 3554 32450 3566
rect 32398 3490 32450 3502
rect 35310 3554 35362 3566
rect 35310 3490 35362 3502
rect 39118 3554 39170 3566
rect 39118 3490 39170 3502
rect 39566 3554 39618 3566
rect 39566 3490 39618 3502
rect 39790 3554 39842 3566
rect 39790 3490 39842 3502
rect 40910 3554 40962 3566
rect 40910 3490 40962 3502
rect 41358 3554 41410 3566
rect 41358 3490 41410 3502
rect 41582 3554 41634 3566
rect 41582 3490 41634 3502
rect 39342 3442 39394 3454
rect 3826 3390 3838 3442
rect 3890 3390 3902 3442
rect 8754 3390 8766 3442
rect 8818 3390 8830 3442
rect 22530 3390 22542 3442
rect 22594 3390 22606 3442
rect 26338 3390 26350 3442
rect 26402 3390 26414 3442
rect 30258 3390 30270 3442
rect 30322 3390 30334 3442
rect 34514 3390 34526 3442
rect 34578 3390 34590 3442
rect 38098 3390 38110 3442
rect 38162 3390 38174 3442
rect 39342 3378 39394 3390
rect 41470 3442 41522 3454
rect 41470 3378 41522 3390
rect 32510 3330 32562 3342
rect 32510 3266 32562 3278
rect 35422 3330 35474 3342
rect 35422 3266 35474 3278
rect 40126 3330 40178 3342
rect 40126 3266 40178 3278
rect 1344 3162 42560 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 42560 3162
rect 1344 3076 42560 3110
<< via1 >>
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 30158 24558 30210 24610
rect 30606 24558 30658 24610
rect 31838 24558 31890 24610
rect 41582 24558 41634 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 32062 24110 32114 24162
rect 32958 24110 33010 24162
rect 28030 23998 28082 24050
rect 30494 23998 30546 24050
rect 32958 23998 33010 24050
rect 35758 23998 35810 24050
rect 36878 23998 36930 24050
rect 34190 23886 34242 23938
rect 39454 23774 39506 23826
rect 28702 23662 28754 23714
rect 29598 23662 29650 23714
rect 30046 23662 30098 23714
rect 31166 23662 31218 23714
rect 31502 23662 31554 23714
rect 32062 23662 32114 23714
rect 32510 23662 32562 23714
rect 33294 23662 33346 23714
rect 33854 23662 33906 23714
rect 35310 23662 35362 23714
rect 36430 23662 36482 23714
rect 37774 23662 37826 23714
rect 38222 23662 38274 23714
rect 38670 23662 38722 23714
rect 39118 23662 39170 23714
rect 40238 23662 40290 23714
rect 40686 23662 40738 23714
rect 41358 23662 41410 23714
rect 41806 23662 41858 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 32958 23326 33010 23378
rect 32510 23214 32562 23266
rect 39678 23214 39730 23266
rect 42030 23214 42082 23266
rect 29710 23102 29762 23154
rect 37662 23102 37714 23154
rect 26238 22990 26290 23042
rect 26574 22990 26626 23042
rect 27134 22990 27186 23042
rect 27582 22990 27634 23042
rect 28254 22990 28306 23042
rect 28590 22990 28642 23042
rect 29374 22990 29426 23042
rect 30494 22990 30546 23042
rect 30830 22990 30882 23042
rect 31614 22990 31666 23042
rect 31950 22990 32002 23042
rect 33518 22990 33570 23042
rect 33966 22990 34018 23042
rect 34526 22990 34578 23042
rect 34862 22990 34914 23042
rect 35422 22990 35474 23042
rect 35870 22990 35922 23042
rect 36206 22990 36258 23042
rect 36766 22990 36818 23042
rect 37102 22990 37154 23042
rect 38334 22990 38386 23042
rect 38782 22990 38834 23042
rect 39230 22990 39282 23042
rect 40238 22990 40290 23042
rect 40686 22990 40738 23042
rect 41470 22990 41522 23042
rect 35646 22878 35698 22930
rect 36766 22878 36818 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 35982 22542 36034 22594
rect 36430 22542 36482 22594
rect 3278 22430 3330 22482
rect 24782 22430 24834 22482
rect 25230 22430 25282 22482
rect 25566 22430 25618 22482
rect 26014 22430 26066 22482
rect 26462 22430 26514 22482
rect 29486 22430 29538 22482
rect 30046 22430 30098 22482
rect 31390 22430 31442 22482
rect 31726 22430 31778 22482
rect 32174 22430 32226 22482
rect 32622 22430 32674 22482
rect 34190 22430 34242 22482
rect 35086 22430 35138 22482
rect 36430 22430 36482 22482
rect 38558 22430 38610 22482
rect 38894 22430 38946 22482
rect 30494 22318 30546 22370
rect 37886 22318 37938 22370
rect 38894 22318 38946 22370
rect 1934 22206 1986 22258
rect 27806 22206 27858 22258
rect 38334 22206 38386 22258
rect 40014 22206 40066 22258
rect 26910 22094 26962 22146
rect 27470 22094 27522 22146
rect 28590 22094 28642 22146
rect 30942 22094 30994 22146
rect 33406 22094 33458 22146
rect 33742 22094 33794 22146
rect 34750 22094 34802 22146
rect 35534 22094 35586 22146
rect 35982 22094 36034 22146
rect 37438 22094 37490 22146
rect 40574 22094 40626 22146
rect 41022 22094 41074 22146
rect 41694 22094 41746 22146
rect 42030 22094 42082 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 1822 21758 1874 21810
rect 28814 21758 28866 21810
rect 32174 21758 32226 21810
rect 34862 21758 34914 21810
rect 35758 21758 35810 21810
rect 37550 21758 37602 21810
rect 38894 21758 38946 21810
rect 42030 21758 42082 21810
rect 26686 21534 26738 21586
rect 34078 21534 34130 21586
rect 24110 21422 24162 21474
rect 24558 21422 24610 21474
rect 24894 21422 24946 21474
rect 25566 21422 25618 21474
rect 26238 21422 26290 21474
rect 27134 21422 27186 21474
rect 27582 21422 27634 21474
rect 28030 21422 28082 21474
rect 28478 21422 28530 21474
rect 29262 21422 29314 21474
rect 30158 21422 30210 21474
rect 30494 21422 30546 21474
rect 31054 21422 31106 21474
rect 31726 21422 31778 21474
rect 32734 21422 32786 21474
rect 33630 21422 33682 21474
rect 34414 21422 34466 21474
rect 35422 21422 35474 21474
rect 36318 21422 36370 21474
rect 36766 21422 36818 21474
rect 37214 21422 37266 21474
rect 37998 21422 38050 21474
rect 38446 21422 38498 21474
rect 39342 21422 39394 21474
rect 40014 21422 40066 21474
rect 40462 21422 40514 21474
rect 41470 21422 41522 21474
rect 37214 21310 37266 21362
rect 38110 21310 38162 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 33518 20974 33570 21026
rect 34414 20974 34466 21026
rect 34862 20974 34914 21026
rect 35086 20974 35138 21026
rect 35310 20974 35362 21026
rect 36206 20974 36258 21026
rect 22990 20862 23042 20914
rect 23438 20862 23490 20914
rect 23886 20862 23938 20914
rect 29934 20862 29986 20914
rect 31278 20862 31330 20914
rect 32622 20862 32674 20914
rect 33070 20862 33122 20914
rect 33518 20862 33570 20914
rect 34414 20862 34466 20914
rect 34862 20862 34914 20914
rect 35310 20862 35362 20914
rect 35758 20862 35810 20914
rect 38782 20862 38834 20914
rect 41246 20862 41298 20914
rect 42030 20862 42082 20914
rect 26238 20750 26290 20802
rect 36206 20750 36258 20802
rect 37438 20750 37490 20802
rect 24334 20638 24386 20690
rect 26574 20638 26626 20690
rect 28702 20638 28754 20690
rect 36654 20638 36706 20690
rect 24670 20526 24722 20578
rect 25230 20526 25282 20578
rect 25790 20526 25842 20578
rect 27022 20526 27074 20578
rect 27918 20526 27970 20578
rect 28366 20526 28418 20578
rect 29486 20526 29538 20578
rect 30494 20526 30546 20578
rect 30942 20526 30994 20578
rect 31838 20526 31890 20578
rect 32286 20526 32338 20578
rect 33966 20526 34018 20578
rect 37886 20526 37938 20578
rect 38334 20526 38386 20578
rect 39230 20526 39282 20578
rect 40014 20526 40066 20578
rect 40462 20526 40514 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 31838 20190 31890 20242
rect 34862 20190 34914 20242
rect 22878 20078 22930 20130
rect 23326 20078 23378 20130
rect 25566 20078 25618 20130
rect 39342 20078 39394 20130
rect 26014 19966 26066 20018
rect 27806 19966 27858 20018
rect 33518 19966 33570 20018
rect 34414 19966 34466 20018
rect 37998 19966 38050 20018
rect 22094 19854 22146 19906
rect 22542 19854 22594 19906
rect 23886 19854 23938 19906
rect 24222 19854 24274 19906
rect 24670 19854 24722 19906
rect 26574 19854 26626 19906
rect 26910 19854 26962 19906
rect 27470 19854 27522 19906
rect 28254 19854 28306 19906
rect 28702 19854 28754 19906
rect 29262 19854 29314 19906
rect 29598 19854 29650 19906
rect 30158 19854 30210 19906
rect 30494 19854 30546 19906
rect 31054 19854 31106 19906
rect 31390 19854 31442 19906
rect 32286 19854 32338 19906
rect 32846 19854 32898 19906
rect 33966 19854 34018 19906
rect 35422 19854 35474 19906
rect 35758 19854 35810 19906
rect 36206 19854 36258 19906
rect 36766 19854 36818 19906
rect 37102 19854 37154 19906
rect 37550 19854 37602 19906
rect 38446 19854 38498 19906
rect 38894 19854 38946 19906
rect 39790 19854 39842 19906
rect 40350 19854 40402 19906
rect 40798 19854 40850 19906
rect 41470 19854 41522 19906
rect 41918 19854 41970 19906
rect 21982 19742 22034 19794
rect 23326 19742 23378 19794
rect 28702 19742 28754 19794
rect 29486 19742 29538 19794
rect 37326 19742 37378 19794
rect 37886 19742 37938 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 37438 19406 37490 19458
rect 38334 19406 38386 19458
rect 39678 19406 39730 19458
rect 40238 19406 40290 19458
rect 41246 19406 41298 19458
rect 41918 19406 41970 19458
rect 21646 19294 21698 19346
rect 27694 19294 27746 19346
rect 28590 19294 28642 19346
rect 33630 19294 33682 19346
rect 35086 19294 35138 19346
rect 37886 19294 37938 19346
rect 40238 19294 40290 19346
rect 42030 19294 42082 19346
rect 23326 19182 23378 19234
rect 23662 19182 23714 19234
rect 25230 19182 25282 19234
rect 34190 19182 34242 19234
rect 25006 19070 25058 19122
rect 25902 19070 25954 19122
rect 26238 19070 26290 19122
rect 39678 19070 39730 19122
rect 20862 18958 20914 19010
rect 22094 18958 22146 19010
rect 22542 18958 22594 19010
rect 22990 18958 23042 19010
rect 23550 18958 23602 19010
rect 24110 18958 24162 19010
rect 25454 18958 25506 19010
rect 25566 18958 25618 19010
rect 26126 18958 26178 19010
rect 26686 18958 26738 19010
rect 27134 18958 27186 19010
rect 28142 18958 28194 19010
rect 29486 18958 29538 19010
rect 29934 18958 29986 19010
rect 30718 18958 30770 19010
rect 31166 18958 31218 19010
rect 31614 18958 31666 19010
rect 32286 18958 32338 19010
rect 32846 18958 32898 19010
rect 33294 18958 33346 19010
rect 34638 18958 34690 19010
rect 35758 18958 35810 19010
rect 36206 18958 36258 19010
rect 36654 18958 36706 19010
rect 37438 18958 37490 19010
rect 38334 18958 38386 19010
rect 38782 18958 38834 19010
rect 39230 18958 39282 19010
rect 40686 18958 40738 19010
rect 41246 18958 41298 19010
rect 41694 18958 41746 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 24110 18622 24162 18674
rect 29822 18622 29874 18674
rect 24334 18510 24386 18562
rect 20638 18398 20690 18450
rect 23886 18398 23938 18450
rect 24446 18398 24498 18450
rect 26126 18398 26178 18450
rect 29934 18398 29986 18450
rect 36094 18398 36146 18450
rect 36318 18398 36370 18450
rect 39006 18398 39058 18450
rect 39454 18398 39506 18450
rect 41918 18398 41970 18450
rect 20078 18286 20130 18338
rect 21310 18286 21362 18338
rect 23438 18286 23490 18338
rect 26798 18286 26850 18338
rect 28926 18286 28978 18338
rect 30606 18286 30658 18338
rect 31054 18286 31106 18338
rect 31502 18286 31554 18338
rect 31950 18286 32002 18338
rect 32398 18286 32450 18338
rect 32958 18286 33010 18338
rect 33518 18286 33570 18338
rect 34078 18286 34130 18338
rect 34862 18286 34914 18338
rect 35422 18286 35474 18338
rect 35870 18286 35922 18338
rect 36430 18286 36482 18338
rect 37102 18286 37154 18338
rect 37662 18286 37714 18338
rect 38110 18286 38162 18338
rect 38558 18286 38610 18338
rect 39902 18286 39954 18338
rect 40462 18286 40514 18338
rect 40798 18286 40850 18338
rect 42030 18286 42082 18338
rect 29822 18174 29874 18226
rect 30494 18174 30546 18226
rect 34974 18174 35026 18226
rect 35534 18174 35586 18226
rect 35870 18174 35922 18226
rect 36542 18174 36594 18226
rect 37214 18174 37266 18226
rect 37886 18174 37938 18226
rect 38558 18174 38610 18226
rect 40350 18174 40402 18226
rect 40798 18174 40850 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 23438 17838 23490 17890
rect 24782 17838 24834 17890
rect 25454 17838 25506 17890
rect 25790 17838 25842 17890
rect 27358 17838 27410 17890
rect 28142 17838 28194 17890
rect 41246 17838 41298 17890
rect 42030 17838 42082 17890
rect 18622 17726 18674 17778
rect 19070 17726 19122 17778
rect 19854 17726 19906 17778
rect 20862 17726 20914 17778
rect 21758 17726 21810 17778
rect 26014 17726 26066 17778
rect 28590 17726 28642 17778
rect 30942 17726 30994 17778
rect 35310 17726 35362 17778
rect 41358 17726 41410 17778
rect 41918 17726 41970 17778
rect 21646 17614 21698 17666
rect 21870 17614 21922 17666
rect 22318 17614 22370 17666
rect 23774 17614 23826 17666
rect 24110 17614 24162 17666
rect 30046 17614 30098 17666
rect 30270 17614 30322 17666
rect 32510 17614 32562 17666
rect 38782 17614 38834 17666
rect 23550 17502 23602 17554
rect 24894 17502 24946 17554
rect 26574 17502 26626 17554
rect 26910 17502 26962 17554
rect 27470 17502 27522 17554
rect 28030 17502 28082 17554
rect 31054 17502 31106 17554
rect 33182 17502 33234 17554
rect 35982 17502 36034 17554
rect 37550 17502 37602 17554
rect 39230 17502 39282 17554
rect 40574 17502 40626 17554
rect 19518 17390 19570 17442
rect 20414 17390 20466 17442
rect 22990 17390 23042 17442
rect 24782 17390 24834 17442
rect 26686 17390 26738 17442
rect 29822 17390 29874 17442
rect 30158 17390 30210 17442
rect 30830 17390 30882 17442
rect 31278 17390 31330 17442
rect 31838 17390 31890 17442
rect 36094 17390 36146 17442
rect 36318 17390 36370 17442
rect 36654 17390 36706 17442
rect 37662 17390 37714 17442
rect 38110 17390 38162 17442
rect 38222 17390 38274 17442
rect 38446 17390 38498 17442
rect 39342 17390 39394 17442
rect 40014 17390 40066 17442
rect 40686 17390 40738 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 18734 17054 18786 17106
rect 19518 17054 19570 17106
rect 19966 17054 20018 17106
rect 21310 17054 21362 17106
rect 23102 17054 23154 17106
rect 24446 17054 24498 17106
rect 26238 17054 26290 17106
rect 31614 17054 31666 17106
rect 32174 17054 32226 17106
rect 37102 17054 37154 17106
rect 37326 17054 37378 17106
rect 38670 17054 38722 17106
rect 21758 16942 21810 16994
rect 23326 16942 23378 16994
rect 23438 16942 23490 16994
rect 24222 16942 24274 16994
rect 30942 16942 30994 16994
rect 31390 16942 31442 16994
rect 31726 16942 31778 16994
rect 32398 16942 32450 16994
rect 38334 16942 38386 16994
rect 39566 16942 39618 16994
rect 40574 16942 40626 16994
rect 41806 16942 41858 16994
rect 41918 16942 41970 16994
rect 15262 16830 15314 16882
rect 17614 16830 17666 16882
rect 18286 16830 18338 16882
rect 20414 16830 20466 16882
rect 20862 16830 20914 16882
rect 22206 16830 22258 16882
rect 22654 16830 22706 16882
rect 24110 16830 24162 16882
rect 24894 16830 24946 16882
rect 27022 16830 27074 16882
rect 30382 16830 30434 16882
rect 30718 16830 30770 16882
rect 32510 16830 32562 16882
rect 33630 16830 33682 16882
rect 34414 16830 34466 16882
rect 37662 16830 37714 16882
rect 38558 16830 38610 16882
rect 39006 16830 39058 16882
rect 39342 16830 39394 16882
rect 39678 16830 39730 16882
rect 40462 16830 40514 16882
rect 19070 16718 19122 16770
rect 25678 16718 25730 16770
rect 27806 16718 27858 16770
rect 29934 16718 29986 16770
rect 30830 16718 30882 16770
rect 36542 16718 36594 16770
rect 37214 16718 37266 16770
rect 25902 16606 25954 16658
rect 41806 16606 41858 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15374 16270 15426 16322
rect 16270 16270 16322 16322
rect 20414 16270 20466 16322
rect 20750 16270 20802 16322
rect 14366 16158 14418 16210
rect 16270 16158 16322 16210
rect 18734 16158 18786 16210
rect 19182 16158 19234 16210
rect 20414 16158 20466 16210
rect 23214 16158 23266 16210
rect 24670 16158 24722 16210
rect 21982 16046 22034 16098
rect 22318 16046 22370 16098
rect 22990 16046 23042 16098
rect 24110 16046 24162 16098
rect 24334 16046 24386 16098
rect 25454 16046 25506 16098
rect 25902 16046 25954 16098
rect 21646 15934 21698 15986
rect 23102 15934 23154 15986
rect 25230 15934 25282 15986
rect 26014 15934 26066 15986
rect 26798 16270 26850 16322
rect 33854 16270 33906 16322
rect 39902 16270 39954 16322
rect 26350 16158 26402 16210
rect 27358 16158 27410 16210
rect 28366 16158 28418 16210
rect 30718 16158 30770 16210
rect 33182 16158 33234 16210
rect 37662 16158 37714 16210
rect 38782 16158 38834 16210
rect 39566 16158 39618 16210
rect 27022 16046 27074 16098
rect 27246 16046 27298 16098
rect 27470 16046 27522 16098
rect 28030 16046 28082 16098
rect 28254 16046 28306 16098
rect 28702 16046 28754 16098
rect 30158 16046 30210 16098
rect 31278 16046 31330 16098
rect 31838 16046 31890 16098
rect 32846 16046 32898 16098
rect 33070 16046 33122 16098
rect 33294 16046 33346 16098
rect 35310 16046 35362 16098
rect 35646 16046 35698 16098
rect 35982 16046 36034 16098
rect 36318 16046 36370 16098
rect 37438 16046 37490 16098
rect 39118 16046 39170 16098
rect 41806 16046 41858 16098
rect 31502 15934 31554 15986
rect 32622 15934 32674 15986
rect 33966 15934 34018 15986
rect 34638 15934 34690 15986
rect 34750 15934 34802 15986
rect 35422 15934 35474 15986
rect 36542 15934 36594 15986
rect 37998 15934 38050 15986
rect 38782 15934 38834 15986
rect 39790 15934 39842 15986
rect 40574 15934 40626 15986
rect 41694 15934 41746 15986
rect 14926 15822 14978 15874
rect 15374 15822 15426 15874
rect 15710 15822 15762 15874
rect 16718 15822 16770 15874
rect 17166 15822 17218 15874
rect 17614 15822 17666 15874
rect 17950 15822 18002 15874
rect 19742 15822 19794 15874
rect 20862 15822 20914 15874
rect 21982 15822 22034 15874
rect 23326 15822 23378 15874
rect 23438 15822 23490 15874
rect 25566 15822 25618 15874
rect 25678 15822 25730 15874
rect 28478 15822 28530 15874
rect 29486 15822 29538 15874
rect 29598 15822 29650 15874
rect 29822 15822 29874 15874
rect 30606 15822 30658 15874
rect 31390 15822 31442 15874
rect 34414 15822 34466 15874
rect 36654 15822 36706 15874
rect 37774 15822 37826 15874
rect 38558 15822 38610 15874
rect 40462 15822 40514 15874
rect 41022 15822 41074 15874
rect 41470 15822 41522 15874
rect 42030 15822 42082 15874
rect 42254 15822 42306 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 13358 15486 13410 15538
rect 14590 15486 14642 15538
rect 18286 15486 18338 15538
rect 19966 15486 20018 15538
rect 23886 15486 23938 15538
rect 24110 15486 24162 15538
rect 25902 15486 25954 15538
rect 26910 15486 26962 15538
rect 27134 15486 27186 15538
rect 30382 15486 30434 15538
rect 30606 15486 30658 15538
rect 31502 15486 31554 15538
rect 31614 15486 31666 15538
rect 35646 15486 35698 15538
rect 35870 15486 35922 15538
rect 36430 15486 36482 15538
rect 36654 15486 36706 15538
rect 37214 15486 37266 15538
rect 39790 15486 39842 15538
rect 40574 15486 40626 15538
rect 41806 15486 41858 15538
rect 42030 15486 42082 15538
rect 21310 15374 21362 15426
rect 24222 15374 24274 15426
rect 24670 15374 24722 15426
rect 26238 15374 26290 15426
rect 28702 15374 28754 15426
rect 29486 15374 29538 15426
rect 29934 15374 29986 15426
rect 31726 15374 31778 15426
rect 32398 15374 32450 15426
rect 33742 15374 33794 15426
rect 33854 15374 33906 15426
rect 36318 15374 36370 15426
rect 37102 15374 37154 15426
rect 37438 15374 37490 15426
rect 38334 15374 38386 15426
rect 39454 15374 39506 15426
rect 39566 15374 39618 15426
rect 40350 15374 40402 15426
rect 20638 15262 20690 15314
rect 25566 15262 25618 15314
rect 26014 15262 26066 15314
rect 26798 15262 26850 15314
rect 27470 15262 27522 15314
rect 28142 15262 28194 15314
rect 28478 15262 28530 15314
rect 29374 15262 29426 15314
rect 29710 15262 29762 15314
rect 30718 15262 30770 15314
rect 32286 15262 32338 15314
rect 33518 15262 33570 15314
rect 34974 15262 35026 15314
rect 35534 15262 35586 15314
rect 38670 15262 38722 15314
rect 38782 15262 38834 15314
rect 38894 15262 38946 15314
rect 40238 15262 40290 15314
rect 41694 15318 41746 15370
rect 11678 15150 11730 15202
rect 12574 15150 12626 15202
rect 13022 15150 13074 15202
rect 13918 15150 13970 15202
rect 15262 15150 15314 15202
rect 15822 15150 15874 15202
rect 16494 15150 16546 15202
rect 16942 15150 16994 15202
rect 17838 15150 17890 15202
rect 18846 15150 18898 15202
rect 19182 15150 19234 15202
rect 23438 15150 23490 15202
rect 28814 15150 28866 15202
rect 34862 15150 34914 15202
rect 37774 15150 37826 15202
rect 24446 15038 24498 15090
rect 25118 15038 25170 15090
rect 32398 15038 32450 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 11230 14702 11282 14754
rect 11678 14702 11730 14754
rect 16942 14702 16994 14754
rect 17278 14702 17330 14754
rect 27246 14702 27298 14754
rect 31278 14702 31330 14754
rect 34190 14702 34242 14754
rect 9662 14590 9714 14642
rect 10110 14590 10162 14642
rect 18622 14590 18674 14642
rect 24558 14590 24610 14642
rect 25118 14590 25170 14642
rect 27918 14590 27970 14642
rect 32734 14590 32786 14642
rect 34862 14590 34914 14642
rect 36206 14590 36258 14642
rect 20078 14478 20130 14530
rect 21758 14478 21810 14530
rect 27134 14478 27186 14530
rect 29598 14478 29650 14530
rect 30270 14478 30322 14530
rect 31390 14478 31442 14530
rect 32398 14478 32450 14530
rect 32622 14478 32674 14530
rect 32846 14478 32898 14530
rect 33294 14478 33346 14530
rect 33630 14478 33682 14530
rect 38782 14478 38834 14530
rect 40350 14478 40402 14530
rect 41806 14478 41858 14530
rect 20190 14366 20242 14418
rect 22430 14366 22482 14418
rect 26462 14366 26514 14418
rect 28814 14366 28866 14418
rect 29710 14366 29762 14418
rect 30606 14366 30658 14418
rect 32174 14366 32226 14418
rect 33518 14366 33570 14418
rect 34302 14366 34354 14418
rect 36094 14366 36146 14418
rect 37662 14366 37714 14418
rect 39118 14366 39170 14418
rect 39566 14366 39618 14418
rect 39902 14366 39954 14418
rect 40686 14366 40738 14418
rect 9214 14254 9266 14306
rect 11118 14254 11170 14306
rect 11566 14254 11618 14306
rect 11902 14254 11954 14306
rect 12462 14254 12514 14306
rect 12910 14254 12962 14306
rect 13582 14254 13634 14306
rect 14142 14254 14194 14306
rect 14478 14254 14530 14306
rect 15038 14254 15090 14306
rect 15598 14254 15650 14306
rect 16046 14254 16098 14306
rect 16494 14254 16546 14306
rect 16942 14254 16994 14306
rect 17390 14254 17442 14306
rect 18174 14254 18226 14306
rect 19070 14254 19122 14306
rect 19630 14254 19682 14306
rect 20414 14254 20466 14306
rect 20862 14254 20914 14306
rect 25230 14254 25282 14306
rect 25902 14254 25954 14306
rect 26574 14254 26626 14306
rect 27246 14254 27298 14306
rect 28590 14254 28642 14306
rect 28702 14254 28754 14306
rect 29934 14254 29986 14306
rect 30494 14254 30546 14306
rect 31278 14254 31330 14306
rect 34974 14254 35026 14306
rect 35422 14254 35474 14306
rect 36318 14254 36370 14306
rect 36542 14254 36594 14306
rect 37550 14254 37602 14306
rect 38110 14254 38162 14306
rect 38894 14254 38946 14306
rect 40574 14254 40626 14306
rect 41470 14254 41522 14306
rect 41694 14254 41746 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 15150 13918 15202 13970
rect 15598 13918 15650 13970
rect 16606 13918 16658 13970
rect 16942 13918 16994 13970
rect 24110 13918 24162 13970
rect 27022 13918 27074 13970
rect 32734 13918 32786 13970
rect 33854 13918 33906 13970
rect 34862 13918 34914 13970
rect 36206 13918 36258 13970
rect 36654 13918 36706 13970
rect 39454 13918 39506 13970
rect 39566 13918 39618 13970
rect 40014 13918 40066 13970
rect 41694 13918 41746 13970
rect 14254 13806 14306 13858
rect 21310 13806 21362 13858
rect 21534 13806 21586 13858
rect 21646 13806 21698 13858
rect 22766 13806 22818 13858
rect 24782 13806 24834 13858
rect 28478 13806 28530 13858
rect 32510 13806 32562 13858
rect 32846 13806 32898 13858
rect 33630 13806 33682 13858
rect 35982 13806 36034 13858
rect 37214 13806 37266 13858
rect 38334 13806 38386 13858
rect 40686 13806 40738 13858
rect 13358 13694 13410 13746
rect 17950 13694 18002 13746
rect 21982 13694 22034 13746
rect 22878 13694 22930 13746
rect 24894 13694 24946 13746
rect 25678 13694 25730 13746
rect 25902 13694 25954 13746
rect 26350 13694 26402 13746
rect 26798 13694 26850 13746
rect 26910 13694 26962 13746
rect 27358 13694 27410 13746
rect 28030 13694 28082 13746
rect 29262 13694 29314 13746
rect 34078 13694 34130 13746
rect 34302 13694 34354 13746
rect 35870 13694 35922 13746
rect 38894 13694 38946 13746
rect 39342 13694 39394 13746
rect 40574 13694 40626 13746
rect 40910 13694 40962 13746
rect 41582 13694 41634 13746
rect 6750 13582 6802 13634
rect 7198 13582 7250 13634
rect 7646 13582 7698 13634
rect 8094 13582 8146 13634
rect 8654 13582 8706 13634
rect 8990 13582 9042 13634
rect 9886 13582 9938 13634
rect 10334 13582 10386 13634
rect 11118 13582 11170 13634
rect 11678 13582 11730 13634
rect 12014 13582 12066 13634
rect 12574 13582 12626 13634
rect 12910 13582 12962 13634
rect 13918 13582 13970 13634
rect 14702 13582 14754 13634
rect 16046 13582 16098 13634
rect 18622 13582 18674 13634
rect 20750 13582 20802 13634
rect 22094 13582 22146 13634
rect 23550 13582 23602 13634
rect 25790 13582 25842 13634
rect 29934 13582 29986 13634
rect 32062 13582 32114 13634
rect 33966 13582 34018 13634
rect 34974 13582 35026 13634
rect 38446 13582 38498 13634
rect 6750 13470 6802 13522
rect 7422 13470 7474 13522
rect 7646 13470 7698 13522
rect 8878 13470 8930 13522
rect 9214 13470 9266 13522
rect 12574 13470 12626 13522
rect 13246 13470 13298 13522
rect 13582 13470 13634 13522
rect 14142 13470 14194 13522
rect 16158 13470 16210 13522
rect 16606 13470 16658 13522
rect 22766 13470 22818 13522
rect 24782 13470 24834 13522
rect 36990 13470 37042 13522
rect 38110 13470 38162 13522
rect 41694 13470 41746 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 27806 13134 27858 13186
rect 36654 13134 36706 13186
rect 6414 13022 6466 13074
rect 7198 13022 7250 13074
rect 12686 13022 12738 13074
rect 20414 13022 20466 13074
rect 22990 13022 23042 13074
rect 27134 13022 27186 13074
rect 29710 13022 29762 13074
rect 33070 13022 33122 13074
rect 35198 13022 35250 13074
rect 37774 13022 37826 13074
rect 10110 12910 10162 12962
rect 12126 12910 12178 12962
rect 13694 12910 13746 12962
rect 19070 12910 19122 12962
rect 19742 12910 19794 12962
rect 20750 12910 20802 12962
rect 23438 12910 23490 12962
rect 24222 12910 24274 12962
rect 29486 12910 29538 12962
rect 30158 12910 30210 12962
rect 31054 12910 31106 12962
rect 32398 12910 32450 12962
rect 35758 12910 35810 12962
rect 38222 12910 38274 12962
rect 38670 12910 38722 12962
rect 39342 12910 39394 12962
rect 39678 12910 39730 12962
rect 40014 12910 40066 12962
rect 40574 12910 40626 12962
rect 41470 12910 41522 12962
rect 41806 12910 41858 12962
rect 9326 12798 9378 12850
rect 10782 12798 10834 12850
rect 12014 12798 12066 12850
rect 12798 12798 12850 12850
rect 12910 12798 12962 12850
rect 13134 12798 13186 12850
rect 14478 12798 14530 12850
rect 17278 12798 17330 12850
rect 17838 12798 17890 12850
rect 18510 12798 18562 12850
rect 21982 12798 22034 12850
rect 25006 12798 25058 12850
rect 27694 12798 27746 12850
rect 28366 12798 28418 12850
rect 29934 12798 29986 12850
rect 30718 12798 30770 12850
rect 30830 12798 30882 12850
rect 31502 12798 31554 12850
rect 31614 12798 31666 12850
rect 35870 12798 35922 12850
rect 36094 12798 36146 12850
rect 36654 12798 36706 12850
rect 36766 12798 36818 12850
rect 37662 12798 37714 12850
rect 37998 12798 38050 12850
rect 39006 12798 39058 12850
rect 39902 12798 39954 12850
rect 5966 12686 6018 12738
rect 10670 12686 10722 12738
rect 11454 12686 11506 12738
rect 13806 12686 13858 12738
rect 14030 12686 14082 12738
rect 14590 12686 14642 12738
rect 15486 12686 15538 12738
rect 15934 12686 15986 12738
rect 16270 12686 16322 12738
rect 16830 12686 16882 12738
rect 17726 12686 17778 12738
rect 18398 12686 18450 12738
rect 19406 12686 19458 12738
rect 19630 12686 19682 12738
rect 22094 12686 22146 12738
rect 22878 12686 22930 12738
rect 23102 12686 23154 12738
rect 27918 12686 27970 12738
rect 28142 12686 28194 12738
rect 28814 12686 28866 12738
rect 31838 12686 31890 12738
rect 38782 12686 38834 12738
rect 40686 12686 40738 12738
rect 40910 12686 40962 12738
rect 41694 12686 41746 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 12798 12350 12850 12402
rect 15150 12350 15202 12402
rect 15822 12350 15874 12402
rect 16382 12350 16434 12402
rect 29486 12350 29538 12402
rect 30606 12350 30658 12402
rect 32846 12350 32898 12402
rect 33742 12350 33794 12402
rect 35534 12350 35586 12402
rect 36430 12350 36482 12402
rect 36654 12350 36706 12402
rect 37438 12350 37490 12402
rect 38222 12350 38274 12402
rect 38446 12350 38498 12402
rect 39678 12350 39730 12402
rect 41694 12350 41746 12402
rect 9886 12238 9938 12290
rect 11902 12238 11954 12290
rect 13470 12238 13522 12290
rect 13582 12238 13634 12290
rect 14254 12238 14306 12290
rect 14366 12238 14418 12290
rect 15038 12238 15090 12290
rect 18846 12238 18898 12290
rect 18958 12238 19010 12290
rect 25790 12238 25842 12290
rect 25902 12238 25954 12290
rect 27582 12238 27634 12290
rect 28254 12238 28306 12290
rect 28926 12238 28978 12290
rect 29822 12238 29874 12290
rect 33630 12238 33682 12290
rect 34302 12238 34354 12290
rect 34526 12238 34578 12290
rect 35086 12238 35138 12290
rect 36766 12238 36818 12290
rect 37326 12238 37378 12290
rect 38670 12238 38722 12290
rect 39454 12238 39506 12290
rect 40462 12238 40514 12290
rect 40574 12238 40626 12290
rect 41806 12238 41858 12290
rect 6078 12126 6130 12178
rect 10222 12126 10274 12178
rect 11006 12126 11058 12178
rect 12574 12126 12626 12178
rect 12910 12126 12962 12178
rect 14590 12126 14642 12178
rect 15374 12126 15426 12178
rect 19182 12126 19234 12178
rect 23662 12126 23714 12178
rect 25566 12126 25618 12178
rect 26910 12126 26962 12178
rect 27358 12126 27410 12178
rect 28366 12126 28418 12178
rect 29150 12126 29202 12178
rect 29598 12126 29650 12178
rect 30494 12126 30546 12178
rect 30942 12126 30994 12178
rect 31838 12126 31890 12178
rect 33854 12126 33906 12178
rect 35310 12126 35362 12178
rect 35758 12126 35810 12178
rect 36094 12126 36146 12178
rect 4734 12014 4786 12066
rect 5070 12014 5122 12066
rect 5630 12014 5682 12066
rect 6862 12014 6914 12066
rect 8990 12014 9042 12066
rect 11118 12014 11170 12066
rect 12126 12014 12178 12066
rect 16830 12014 16882 12066
rect 17614 12014 17666 12066
rect 18286 12014 18338 12066
rect 21758 12014 21810 12066
rect 30718 12014 30770 12066
rect 32286 12014 32338 12066
rect 39790 12014 39842 12066
rect 9998 11902 10050 11954
rect 10334 11902 10386 11954
rect 11790 11902 11842 11954
rect 13582 11902 13634 11954
rect 16942 11902 16994 11954
rect 17614 11902 17666 11954
rect 17950 11902 18002 11954
rect 18174 11902 18226 11954
rect 26462 11902 26514 11954
rect 27134 11902 27186 11954
rect 28254 11902 28306 11954
rect 29374 11902 29426 11954
rect 31166 11902 31218 11954
rect 34078 11902 34130 11954
rect 35534 11902 35586 11954
rect 37438 11902 37490 11954
rect 38110 11902 38162 11954
rect 40462 11902 40514 11954
rect 41694 11902 41746 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 9662 11566 9714 11618
rect 11006 11566 11058 11618
rect 12798 11566 12850 11618
rect 14814 11566 14866 11618
rect 22542 11566 22594 11618
rect 40462 11566 40514 11618
rect 41918 11566 41970 11618
rect 6862 11454 6914 11506
rect 9886 11454 9938 11506
rect 11790 11454 11842 11506
rect 13918 11454 13970 11506
rect 19406 11454 19458 11506
rect 24222 11454 24274 11506
rect 28702 11454 28754 11506
rect 32174 11454 32226 11506
rect 36766 11454 36818 11506
rect 39454 11454 39506 11506
rect 42030 11454 42082 11506
rect 7086 11342 7138 11394
rect 7758 11342 7810 11394
rect 10894 11342 10946 11394
rect 15934 11342 15986 11394
rect 16606 11342 16658 11394
rect 19966 11342 20018 11394
rect 20190 11342 20242 11394
rect 21870 11342 21922 11394
rect 26910 11342 26962 11394
rect 30158 11342 30210 11394
rect 32846 11342 32898 11394
rect 34638 11342 34690 11394
rect 34862 11342 34914 11394
rect 35086 11342 35138 11394
rect 36094 11342 36146 11394
rect 37774 11342 37826 11394
rect 38222 11342 38274 11394
rect 39790 11342 39842 11394
rect 41358 11342 41410 11394
rect 6078 11230 6130 11282
rect 6750 11230 6802 11282
rect 8094 11230 8146 11282
rect 8654 11230 8706 11282
rect 8990 11230 9042 11282
rect 11678 11230 11730 11282
rect 12126 11230 12178 11282
rect 12910 11230 12962 11282
rect 14142 11230 14194 11282
rect 14702 11230 14754 11282
rect 17278 11230 17330 11282
rect 29598 11230 29650 11282
rect 31390 11230 31442 11282
rect 31950 11230 32002 11282
rect 32958 11230 33010 11282
rect 34190 11230 34242 11282
rect 34414 11230 34466 11282
rect 37662 11230 37714 11282
rect 38446 11230 38498 11282
rect 38558 11230 38610 11282
rect 40462 11230 40514 11282
rect 40574 11230 40626 11282
rect 41246 11230 41298 11282
rect 3614 11118 3666 11170
rect 4062 11118 4114 11170
rect 4510 11118 4562 11170
rect 4958 11118 5010 11170
rect 6190 11118 6242 11170
rect 7646 11118 7698 11170
rect 7870 11118 7922 11170
rect 8878 11118 8930 11170
rect 9886 11118 9938 11170
rect 11006 11118 11058 11170
rect 11902 11118 11954 11170
rect 13918 11118 13970 11170
rect 15374 11118 15426 11170
rect 20526 11118 20578 11170
rect 22206 11118 22258 11170
rect 22430 11118 22482 11170
rect 30046 11118 30098 11170
rect 30830 11118 30882 11170
rect 33182 11118 33234 11170
rect 33518 11118 33570 11170
rect 34526 11118 34578 11170
rect 36094 11118 36146 11170
rect 37438 11118 37490 11170
rect 39566 11118 39618 11170
rect 41022 11118 41074 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 2718 10782 2770 10834
rect 4398 10782 4450 10834
rect 8430 10782 8482 10834
rect 17950 10782 18002 10834
rect 23550 10782 23602 10834
rect 24334 10782 24386 10834
rect 26686 10782 26738 10834
rect 29822 10782 29874 10834
rect 30494 10782 30546 10834
rect 31166 10782 31218 10834
rect 32286 10782 32338 10834
rect 32622 10782 32674 10834
rect 34302 10782 34354 10834
rect 35982 10782 36034 10834
rect 38334 10782 38386 10834
rect 39230 10782 39282 10834
rect 40238 10782 40290 10834
rect 41694 10782 41746 10834
rect 6302 10670 6354 10722
rect 7646 10670 7698 10722
rect 9886 10670 9938 10722
rect 9998 10670 10050 10722
rect 13022 10670 13074 10722
rect 14702 10670 14754 10722
rect 16942 10670 16994 10722
rect 18174 10670 18226 10722
rect 18846 10670 18898 10722
rect 19070 10670 19122 10722
rect 23438 10670 23490 10722
rect 24558 10670 24610 10722
rect 25902 10670 25954 10722
rect 26574 10670 26626 10722
rect 27918 10670 27970 10722
rect 28366 10670 28418 10722
rect 28590 10670 28642 10722
rect 31390 10670 31442 10722
rect 32062 10670 32114 10722
rect 33742 10670 33794 10722
rect 35870 10670 35922 10722
rect 39342 10670 39394 10722
rect 40350 10670 40402 10722
rect 41806 10670 41858 10722
rect 6862 10558 6914 10610
rect 8318 10558 8370 10610
rect 13806 10558 13858 10610
rect 14366 10558 14418 10610
rect 16830 10558 16882 10610
rect 19966 10558 20018 10610
rect 24222 10558 24274 10610
rect 24782 10558 24834 10610
rect 25678 10558 25730 10610
rect 27470 10558 27522 10610
rect 28702 10558 28754 10610
rect 30606 10558 30658 10610
rect 31502 10558 31554 10610
rect 32510 10558 32562 10610
rect 33630 10558 33682 10610
rect 34414 10558 34466 10610
rect 34974 10558 35026 10610
rect 35422 10558 35474 10610
rect 37438 10558 37490 10610
rect 37662 10558 37714 10610
rect 38110 10558 38162 10610
rect 38446 10558 38498 10610
rect 38670 10558 38722 10610
rect 39566 10558 39618 10610
rect 39790 10558 39842 10610
rect 40574 10558 40626 10610
rect 40798 10558 40850 10610
rect 3166 10446 3218 10498
rect 3502 10446 3554 10498
rect 4062 10446 4114 10498
rect 4846 10446 4898 10498
rect 5294 10446 5346 10498
rect 5742 10446 5794 10498
rect 7534 10446 7586 10498
rect 8990 10446 9042 10498
rect 10894 10446 10946 10498
rect 15486 10446 15538 10498
rect 15822 10446 15874 10498
rect 17950 10446 18002 10498
rect 20750 10446 20802 10498
rect 22878 10446 22930 10498
rect 24670 10446 24722 10498
rect 29262 10446 29314 10498
rect 32622 10446 32674 10498
rect 34638 10446 34690 10498
rect 36542 10446 36594 10498
rect 37102 10446 37154 10498
rect 6750 10334 6802 10386
rect 7422 10334 7474 10386
rect 8430 10334 8482 10386
rect 9886 10334 9938 10386
rect 16494 10334 16546 10386
rect 16606 10334 16658 10386
rect 18734 10334 18786 10386
rect 33742 10334 33794 10386
rect 34862 10334 34914 10386
rect 35982 10334 36034 10386
rect 41694 10334 41746 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 2382 9998 2434 10050
rect 3166 9998 3218 10050
rect 10446 9998 10498 10050
rect 12574 9998 12626 10050
rect 17614 9998 17666 10050
rect 19518 9998 19570 10050
rect 21646 9998 21698 10050
rect 30270 9998 30322 10050
rect 36654 9998 36706 10050
rect 37662 9998 37714 10050
rect 2382 9886 2434 9938
rect 2830 9886 2882 9938
rect 4510 9886 4562 9938
rect 5070 9886 5122 9938
rect 6638 9886 6690 9938
rect 10334 9886 10386 9938
rect 13694 9886 13746 9938
rect 19406 9886 19458 9938
rect 20638 9886 20690 9938
rect 20862 9886 20914 9938
rect 22542 9886 22594 9938
rect 24670 9886 24722 9938
rect 25454 9886 25506 9938
rect 27694 9886 27746 9938
rect 30046 9886 30098 9938
rect 30606 9886 30658 9938
rect 33182 9886 33234 9938
rect 35310 9886 35362 9938
rect 36766 9886 36818 9938
rect 38782 9886 38834 9938
rect 39678 9886 39730 9938
rect 9438 9774 9490 9826
rect 11118 9774 11170 9826
rect 11566 9774 11618 9826
rect 11790 9774 11842 9826
rect 16494 9774 16546 9826
rect 17278 9774 17330 9826
rect 17502 9774 17554 9826
rect 18286 9774 18338 9826
rect 19070 9774 19122 9826
rect 19182 9774 19234 9826
rect 21758 9774 21810 9826
rect 22318 9774 22370 9826
rect 22654 9774 22706 9826
rect 23774 9774 23826 9826
rect 26014 9774 26066 9826
rect 26686 9774 26738 9826
rect 27358 9774 27410 9826
rect 28814 9774 28866 9826
rect 31390 9774 31442 9826
rect 31614 9774 31666 9826
rect 32510 9774 32562 9826
rect 37550 9774 37602 9826
rect 37774 9774 37826 9826
rect 38558 9774 38610 9826
rect 39790 9774 39842 9826
rect 40910 9774 40962 9826
rect 6078 9662 6130 9714
rect 8766 9662 8818 9714
rect 12798 9662 12850 9714
rect 15822 9662 15874 9714
rect 17166 9662 17218 9714
rect 21982 9662 22034 9714
rect 23998 9662 24050 9714
rect 24558 9662 24610 9714
rect 25006 9662 25058 9714
rect 27470 9662 27522 9714
rect 27806 9662 27858 9714
rect 31166 9662 31218 9714
rect 35982 9662 36034 9714
rect 36094 9662 36146 9714
rect 37998 9662 38050 9714
rect 39566 9662 39618 9714
rect 40126 9662 40178 9714
rect 40574 9662 40626 9714
rect 40798 9662 40850 9714
rect 41694 9662 41746 9714
rect 1934 9550 1986 9602
rect 3166 9550 3218 9602
rect 3614 9550 3666 9602
rect 4174 9550 4226 9602
rect 5630 9550 5682 9602
rect 10222 9550 10274 9602
rect 11454 9550 11506 9602
rect 12686 9550 12738 9602
rect 18398 9550 18450 9602
rect 18622 9550 18674 9602
rect 23438 9550 23490 9602
rect 23550 9550 23602 9602
rect 24782 9550 24834 9602
rect 26462 9550 26514 9602
rect 26574 9550 26626 9602
rect 28254 9550 28306 9602
rect 28366 9550 28418 9602
rect 28590 9550 28642 9602
rect 29486 9550 29538 9602
rect 31054 9550 31106 9602
rect 35758 9550 35810 9602
rect 38782 9550 38834 9602
rect 41358 9550 41410 9602
rect 41582 9550 41634 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 3838 9214 3890 9266
rect 7982 9214 8034 9266
rect 9886 9214 9938 9266
rect 10894 9214 10946 9266
rect 17726 9214 17778 9266
rect 18286 9214 18338 9266
rect 24558 9214 24610 9266
rect 25566 9214 25618 9266
rect 25678 9214 25730 9266
rect 25902 9214 25954 9266
rect 26910 9214 26962 9266
rect 27134 9214 27186 9266
rect 27246 9214 27298 9266
rect 29710 9214 29762 9266
rect 31054 9214 31106 9266
rect 31278 9214 31330 9266
rect 31838 9214 31890 9266
rect 32062 9214 32114 9266
rect 32734 9214 32786 9266
rect 33854 9214 33906 9266
rect 34638 9214 34690 9266
rect 37326 9214 37378 9266
rect 38110 9214 38162 9266
rect 38894 9214 38946 9266
rect 39454 9214 39506 9266
rect 40462 9214 40514 9266
rect 5406 9102 5458 9154
rect 5966 9102 6018 9154
rect 6078 9102 6130 9154
rect 6862 9102 6914 9154
rect 7086 9102 7138 9154
rect 7534 9102 7586 9154
rect 8878 9102 8930 9154
rect 10110 9102 10162 9154
rect 11902 9102 11954 9154
rect 18510 9102 18562 9154
rect 26126 9102 26178 9154
rect 26686 9102 26738 9154
rect 27806 9102 27858 9154
rect 28590 9102 28642 9154
rect 29038 9102 29090 9154
rect 29598 9102 29650 9154
rect 30830 9102 30882 9154
rect 36654 9102 36706 9154
rect 39678 9102 39730 9154
rect 39790 9102 39842 9154
rect 40574 9102 40626 9154
rect 41694 9102 41746 9154
rect 41806 9102 41858 9154
rect 6302 8990 6354 9042
rect 6750 8990 6802 9042
rect 7758 8990 7810 9042
rect 8206 8990 8258 9042
rect 16718 8990 16770 9042
rect 22430 8990 22482 9042
rect 22990 8990 23042 9042
rect 23438 8990 23490 9042
rect 23550 8990 23602 9042
rect 23662 8990 23714 9042
rect 24110 8990 24162 9042
rect 24782 8990 24834 9042
rect 27918 8990 27970 9042
rect 28478 8990 28530 9042
rect 28814 8990 28866 9042
rect 29934 8990 29986 9042
rect 31390 8990 31442 9042
rect 32286 8990 32338 9042
rect 34750 8990 34802 9042
rect 35422 8990 35474 9042
rect 37438 8990 37490 9042
rect 37998 8990 38050 9042
rect 39006 8990 39058 9042
rect 41470 8990 41522 9042
rect 2158 8878 2210 8930
rect 2494 8878 2546 8930
rect 3054 8878 3106 8930
rect 3390 8878 3442 8930
rect 4286 8878 4338 8930
rect 4734 8878 4786 8930
rect 8990 8878 9042 8930
rect 18174 8878 18226 8930
rect 19182 8878 19234 8930
rect 19630 8878 19682 8930
rect 21758 8878 21810 8930
rect 24670 8878 24722 8930
rect 33966 8878 34018 8930
rect 34862 8878 34914 8930
rect 35534 8878 35586 8930
rect 36318 8878 36370 8930
rect 3390 8766 3442 8818
rect 4510 8766 4562 8818
rect 5294 8766 5346 8818
rect 8654 8766 8706 8818
rect 9774 8766 9826 8818
rect 10670 8766 10722 8818
rect 11006 8766 11058 8818
rect 27806 8766 27858 8818
rect 31726 8766 31778 8818
rect 33630 8766 33682 8818
rect 35758 8766 35810 8818
rect 37326 8766 37378 8818
rect 38110 8766 38162 8818
rect 38894 8766 38946 8818
rect 40462 8766 40514 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 3390 8430 3442 8482
rect 4062 8430 4114 8482
rect 6526 8430 6578 8482
rect 19630 8430 19682 8482
rect 38446 8430 38498 8482
rect 41694 8430 41746 8482
rect 3390 8318 3442 8370
rect 3838 8318 3890 8370
rect 8542 8318 8594 8370
rect 9998 8318 10050 8370
rect 12126 8318 12178 8370
rect 14142 8318 14194 8370
rect 15150 8318 15202 8370
rect 16830 8318 16882 8370
rect 18958 8318 19010 8370
rect 20526 8318 20578 8370
rect 20750 8318 20802 8370
rect 22094 8318 22146 8370
rect 25230 8318 25282 8370
rect 28702 8318 28754 8370
rect 29598 8318 29650 8370
rect 29822 8318 29874 8370
rect 30494 8318 30546 8370
rect 31390 8318 31442 8370
rect 31726 8318 31778 8370
rect 33406 8318 33458 8370
rect 35534 8318 35586 8370
rect 36430 8318 36482 8370
rect 40686 8318 40738 8370
rect 1934 8206 1986 8258
rect 4174 8206 4226 8258
rect 4734 8206 4786 8258
rect 5966 8206 6018 8258
rect 7758 8206 7810 8258
rect 8206 8206 8258 8258
rect 8766 8206 8818 8258
rect 8990 8206 9042 8258
rect 9438 8206 9490 8258
rect 12798 8206 12850 8258
rect 14590 8206 14642 8258
rect 15038 8206 15090 8258
rect 15262 8206 15314 8258
rect 16158 8206 16210 8258
rect 19966 8206 20018 8258
rect 22318 8206 22370 8258
rect 23886 8206 23938 8258
rect 32622 8206 32674 8258
rect 36094 8206 36146 8258
rect 36542 8206 36594 8258
rect 37438 8206 37490 8258
rect 38782 8206 38834 8258
rect 39454 8206 39506 8258
rect 39790 8206 39842 8258
rect 5630 8094 5682 8146
rect 6862 8094 6914 8146
rect 7422 8094 7474 8146
rect 9102 8094 9154 8146
rect 13918 8094 13970 8146
rect 21758 8094 21810 8146
rect 22206 8094 22258 8146
rect 36766 8094 36818 8146
rect 37662 8094 37714 8146
rect 37774 8094 37826 8146
rect 39006 8094 39058 8146
rect 40126 8094 40178 8146
rect 41022 8094 41074 8146
rect 41694 8094 41746 8146
rect 41806 8094 41858 8146
rect 2494 7982 2546 8034
rect 2830 7982 2882 8034
rect 4846 7982 4898 8034
rect 5070 7982 5122 8034
rect 5854 7982 5906 8034
rect 6638 7982 6690 8034
rect 7534 7982 7586 8034
rect 8430 7982 8482 8034
rect 9214 7982 9266 8034
rect 14030 7982 14082 8034
rect 19742 7982 19794 8034
rect 21982 7982 22034 8034
rect 29822 7982 29874 8034
rect 30606 7982 30658 8034
rect 31614 7982 31666 8034
rect 36318 7982 36370 8034
rect 39790 7982 39842 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 1822 7646 1874 7698
rect 2270 7646 2322 7698
rect 2718 7646 2770 7698
rect 3054 7646 3106 7698
rect 6750 7646 6802 7698
rect 7870 7646 7922 7698
rect 8878 7646 8930 7698
rect 10334 7646 10386 7698
rect 10558 7646 10610 7698
rect 21310 7646 21362 7698
rect 23102 7646 23154 7698
rect 25566 7646 25618 7698
rect 26798 7646 26850 7698
rect 29710 7646 29762 7698
rect 30606 7646 30658 7698
rect 31726 7646 31778 7698
rect 33742 7646 33794 7698
rect 35646 7646 35698 7698
rect 36654 7646 36706 7698
rect 37886 7646 37938 7698
rect 37998 7646 38050 7698
rect 38222 7646 38274 7698
rect 39118 7646 39170 7698
rect 40014 7646 40066 7698
rect 41694 7646 41746 7698
rect 3726 7534 3778 7586
rect 4286 7534 4338 7586
rect 4958 7534 5010 7586
rect 5070 7534 5122 7586
rect 5854 7534 5906 7586
rect 6974 7534 7026 7586
rect 10110 7534 10162 7586
rect 21198 7534 21250 7586
rect 21422 7534 21474 7586
rect 22094 7534 22146 7586
rect 22430 7534 22482 7586
rect 23886 7534 23938 7586
rect 26238 7534 26290 7586
rect 27918 7534 27970 7586
rect 32510 7534 32562 7586
rect 35534 7534 35586 7586
rect 36094 7534 36146 7586
rect 39342 7534 39394 7586
rect 39902 7534 39954 7586
rect 41806 7534 41858 7586
rect 4398 7422 4450 7474
rect 5294 7422 5346 7474
rect 5742 7422 5794 7474
rect 6638 7422 6690 7474
rect 7086 7422 7138 7474
rect 8542 7422 8594 7474
rect 8766 7422 8818 7474
rect 8990 7422 9042 7474
rect 10670 7422 10722 7474
rect 16718 7422 16770 7474
rect 17838 7422 17890 7474
rect 22990 7422 23042 7474
rect 23662 7422 23714 7474
rect 26462 7422 26514 7474
rect 27470 7422 27522 7474
rect 28478 7422 28530 7474
rect 28814 7422 28866 7474
rect 29038 7422 29090 7474
rect 30494 7422 30546 7474
rect 30830 7422 30882 7474
rect 31838 7422 31890 7474
rect 32846 7422 32898 7474
rect 34526 7422 34578 7474
rect 34862 7422 34914 7474
rect 36766 7422 36818 7474
rect 36990 7422 37042 7474
rect 38558 7422 38610 7474
rect 40238 7422 40290 7474
rect 3614 7310 3666 7362
rect 6862 7310 6914 7362
rect 7758 7310 7810 7362
rect 11790 7310 11842 7362
rect 18510 7310 18562 7362
rect 20638 7310 20690 7362
rect 23214 7310 23266 7362
rect 24446 7310 24498 7362
rect 24670 7310 24722 7362
rect 28590 7310 28642 7362
rect 29598 7310 29650 7362
rect 31278 7310 31330 7362
rect 32062 7310 32114 7362
rect 33630 7310 33682 7362
rect 35310 7310 35362 7362
rect 36318 7310 36370 7362
rect 37438 7310 37490 7362
rect 39230 7310 39282 7362
rect 40686 7310 40738 7362
rect 5854 7198 5906 7250
rect 10222 7198 10274 7250
rect 23438 7198 23490 7250
rect 29934 7198 29986 7250
rect 32286 7198 32338 7250
rect 33966 7198 34018 7250
rect 35086 7198 35138 7250
rect 36542 7198 36594 7250
rect 41694 7198 41746 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 17278 6862 17330 6914
rect 24110 6862 24162 6914
rect 1934 6750 1986 6802
rect 6526 6750 6578 6802
rect 9998 6750 10050 6802
rect 16830 6750 16882 6802
rect 35086 6750 35138 6802
rect 39006 6750 39058 6802
rect 2382 6638 2434 6690
rect 3278 6638 3330 6690
rect 8654 6638 8706 6690
rect 9438 6638 9490 6690
rect 12798 6638 12850 6690
rect 13918 6638 13970 6690
rect 18622 6638 18674 6690
rect 18958 6638 19010 6690
rect 19406 6638 19458 6690
rect 19854 6638 19906 6690
rect 20638 6638 20690 6690
rect 20974 6638 21026 6690
rect 22766 6638 22818 6690
rect 23214 6638 23266 6690
rect 23438 6638 23490 6690
rect 25454 6638 25506 6690
rect 25678 6638 25730 6690
rect 25902 6638 25954 6690
rect 26350 6638 26402 6690
rect 27022 6638 27074 6690
rect 28142 6638 28194 6690
rect 28702 6638 28754 6690
rect 28814 6638 28866 6690
rect 30158 6638 30210 6690
rect 30382 6638 30434 6690
rect 31390 6638 31442 6690
rect 31614 6638 31666 6690
rect 32286 6638 32338 6690
rect 36654 6638 36706 6690
rect 38446 6638 38498 6690
rect 40910 6638 40962 6690
rect 41582 6638 41634 6690
rect 41918 6638 41970 6690
rect 4174 6526 4226 6578
rect 4846 6526 4898 6578
rect 5966 6526 6018 6578
rect 12126 6526 12178 6578
rect 14702 6526 14754 6578
rect 17390 6526 17442 6578
rect 17838 6526 17890 6578
rect 20078 6526 20130 6578
rect 21646 6526 21698 6578
rect 22206 6526 22258 6578
rect 23998 6526 24050 6578
rect 24670 6526 24722 6578
rect 25230 6526 25282 6578
rect 26798 6526 26850 6578
rect 27694 6526 27746 6578
rect 29710 6526 29762 6578
rect 30942 6526 30994 6578
rect 31278 6526 31330 6578
rect 32958 6526 33010 6578
rect 35982 6526 36034 6578
rect 37886 6526 37938 6578
rect 39902 6526 39954 6578
rect 41022 6526 41074 6578
rect 41806 6526 41858 6578
rect 2718 6414 2770 6466
rect 3726 6414 3778 6466
rect 4286 6414 4338 6466
rect 4958 6414 5010 6466
rect 5630 6414 5682 6466
rect 5854 6414 5906 6466
rect 17614 6414 17666 6466
rect 18398 6414 18450 6466
rect 18510 6414 18562 6466
rect 19630 6414 19682 6466
rect 20750 6414 20802 6466
rect 22990 6414 23042 6466
rect 23102 6414 23154 6466
rect 24222 6414 24274 6466
rect 24446 6414 24498 6466
rect 25566 6414 25618 6466
rect 26686 6414 26738 6466
rect 27918 6414 27970 6466
rect 28030 6414 28082 6466
rect 29934 6414 29986 6466
rect 30046 6414 30098 6466
rect 31166 6414 31218 6466
rect 36206 6414 36258 6466
rect 36318 6414 36370 6466
rect 36430 6414 36482 6466
rect 37774 6414 37826 6466
rect 38110 6414 38162 6466
rect 41246 6414 41298 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 2270 6078 2322 6130
rect 2718 6078 2770 6130
rect 3166 6078 3218 6130
rect 4622 6078 4674 6130
rect 6750 6078 6802 6130
rect 9774 6078 9826 6130
rect 10334 6078 10386 6130
rect 10446 6078 10498 6130
rect 11566 6078 11618 6130
rect 14030 6078 14082 6130
rect 14702 6078 14754 6130
rect 16606 6078 16658 6130
rect 16830 6078 16882 6130
rect 19854 6078 19906 6130
rect 23662 6078 23714 6130
rect 25566 6078 25618 6130
rect 26014 6078 26066 6130
rect 27694 6078 27746 6130
rect 30942 6078 30994 6130
rect 32734 6078 32786 6130
rect 37326 6078 37378 6130
rect 37550 6078 37602 6130
rect 38222 6078 38274 6130
rect 40798 6078 40850 6130
rect 41470 6078 41522 6130
rect 41694 6078 41746 6130
rect 5518 5966 5570 6018
rect 5742 5966 5794 6018
rect 6974 5966 7026 6018
rect 8878 5966 8930 6018
rect 11118 5966 11170 6018
rect 11342 5966 11394 6018
rect 11678 5966 11730 6018
rect 12462 5966 12514 6018
rect 13022 5966 13074 6018
rect 14814 5966 14866 6018
rect 15934 5966 15986 6018
rect 16158 5966 16210 6018
rect 16942 5966 16994 6018
rect 17838 5966 17890 6018
rect 22430 5966 22482 6018
rect 27022 5966 27074 6018
rect 29262 5966 29314 6018
rect 37774 5966 37826 6018
rect 40126 5966 40178 6018
rect 41806 5966 41858 6018
rect 4734 5854 4786 5906
rect 6302 5854 6354 5906
rect 6526 5854 6578 5906
rect 8094 5854 8146 5906
rect 12238 5854 12290 5906
rect 14478 5854 14530 5906
rect 15038 5854 15090 5906
rect 15486 5854 15538 5906
rect 17950 5854 18002 5906
rect 18622 5854 18674 5906
rect 19070 5854 19122 5906
rect 23102 5854 23154 5906
rect 23774 5854 23826 5906
rect 23998 5854 24050 5906
rect 24446 5854 24498 5906
rect 24782 5854 24834 5906
rect 26126 5854 26178 5906
rect 26350 5854 26402 5906
rect 26798 5854 26850 5906
rect 27582 5854 27634 5906
rect 30494 5854 30546 5906
rect 30942 5854 30994 5906
rect 31502 5854 31554 5906
rect 32398 5854 32450 5906
rect 36430 5854 36482 5906
rect 37214 5854 37266 5906
rect 1822 5742 1874 5794
rect 3614 5742 3666 5794
rect 4062 5742 4114 5794
rect 6638 5742 6690 5794
rect 8318 5742 8370 5794
rect 12126 5742 12178 5794
rect 15710 5742 15762 5794
rect 20302 5742 20354 5794
rect 28254 5742 28306 5794
rect 31054 5742 31106 5794
rect 31278 5742 31330 5794
rect 33630 5742 33682 5794
rect 35758 5742 35810 5794
rect 37438 5742 37490 5794
rect 38894 5742 38946 5794
rect 2158 5630 2210 5682
rect 2942 5630 2994 5682
rect 4846 5630 4898 5682
rect 5406 5630 5458 5682
rect 7758 5630 7810 5682
rect 8990 5630 9042 5682
rect 10558 5630 10610 5682
rect 18958 5630 19010 5682
rect 24222 5630 24274 5682
rect 26574 5630 26626 5682
rect 32174 5630 32226 5682
rect 32622 5630 32674 5682
rect 32734 5630 32786 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 3950 5294 4002 5346
rect 6078 5294 6130 5346
rect 23662 5294 23714 5346
rect 24222 5294 24274 5346
rect 25006 5294 25058 5346
rect 28366 5294 28418 5346
rect 35758 5294 35810 5346
rect 35870 5294 35922 5346
rect 41806 5294 41858 5346
rect 2158 5182 2210 5234
rect 2606 5182 2658 5234
rect 3166 5182 3218 5234
rect 6302 5182 6354 5234
rect 6862 5182 6914 5234
rect 8990 5182 9042 5234
rect 10334 5182 10386 5234
rect 12910 5182 12962 5234
rect 13806 5182 13858 5234
rect 15038 5182 15090 5234
rect 17166 5182 17218 5234
rect 18398 5182 18450 5234
rect 20862 5182 20914 5234
rect 22318 5182 22370 5234
rect 25566 5182 25618 5234
rect 28590 5182 28642 5234
rect 31054 5182 31106 5234
rect 31614 5182 31666 5234
rect 33742 5182 33794 5234
rect 37662 5182 37714 5234
rect 39678 5182 39730 5234
rect 4062 5070 4114 5122
rect 5742 5070 5794 5122
rect 9662 5070 9714 5122
rect 12574 5070 12626 5122
rect 14254 5070 14306 5122
rect 17726 5070 17778 5122
rect 19854 5070 19906 5122
rect 21758 5070 21810 5122
rect 23886 5070 23938 5122
rect 24110 5070 24162 5122
rect 27806 5070 27858 5122
rect 28814 5070 28866 5122
rect 36094 5070 36146 5122
rect 36318 5070 36370 5122
rect 41918 5070 41970 5122
rect 4622 4958 4674 5010
rect 10782 4958 10834 5010
rect 11118 4958 11170 5010
rect 11342 4958 11394 5010
rect 11902 4958 11954 5010
rect 12014 4958 12066 5010
rect 19518 4958 19570 5010
rect 19630 4958 19682 5010
rect 20302 4958 20354 5010
rect 24894 4958 24946 5010
rect 26574 4958 26626 5010
rect 28142 4958 28194 5010
rect 29710 4958 29762 5010
rect 32622 4958 32674 5010
rect 34974 4958 35026 5010
rect 38894 4958 38946 5010
rect 40686 4958 40738 5010
rect 41806 4958 41858 5010
rect 3054 4846 3106 4898
rect 3950 4846 4002 4898
rect 4958 4846 5010 4898
rect 10894 4846 10946 4898
rect 12126 4846 12178 4898
rect 23774 4846 23826 4898
rect 28254 4846 28306 4898
rect 36206 4846 36258 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4734 4510 4786 4562
rect 14254 4510 14306 4562
rect 16830 4510 16882 4562
rect 24782 4510 24834 4562
rect 25790 4510 25842 4562
rect 26014 4510 26066 4562
rect 3614 4398 3666 4450
rect 3950 4398 4002 4450
rect 4510 4398 4562 4450
rect 10558 4398 10610 4450
rect 16606 4398 16658 4450
rect 19966 4398 20018 4450
rect 23438 4398 23490 4450
rect 25678 4398 25730 4450
rect 30718 4398 30770 4450
rect 35758 4398 35810 4450
rect 38446 4398 38498 4450
rect 40126 4398 40178 4450
rect 41582 4398 41634 4450
rect 2942 4286 2994 4338
rect 5406 4286 5458 4338
rect 7758 4286 7810 4338
rect 9774 4286 9826 4338
rect 13694 4286 13746 4338
rect 13918 4286 13970 4338
rect 14926 4286 14978 4338
rect 20750 4286 20802 4338
rect 24110 4286 24162 4338
rect 24894 4286 24946 4338
rect 26462 4286 26514 4338
rect 29934 4286 29986 4338
rect 36430 4286 36482 4338
rect 41806 4286 41858 4338
rect 1934 4174 1986 4226
rect 6078 4174 6130 4226
rect 7310 4174 7362 4226
rect 8430 4174 8482 4226
rect 12686 4174 12738 4226
rect 13246 4174 13298 4226
rect 15486 4174 15538 4226
rect 16942 4174 16994 4226
rect 17838 4174 17890 4226
rect 21310 4174 21362 4226
rect 27246 4174 27298 4226
rect 29374 4174 29426 4226
rect 32846 4174 32898 4226
rect 33630 4174 33682 4226
rect 37102 4174 37154 4226
rect 39118 4174 39170 4226
rect 4846 4062 4898 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 21422 3726 21474 3778
rect 31950 3726 32002 3778
rect 35534 3726 35586 3778
rect 35758 3726 35810 3778
rect 2494 3614 2546 3666
rect 6526 3614 6578 3666
rect 10558 3614 10610 3666
rect 12238 3614 12290 3666
rect 14254 3614 14306 3666
rect 16158 3614 16210 3666
rect 18622 3614 18674 3666
rect 20190 3614 20242 3666
rect 21534 3614 21586 3666
rect 24334 3614 24386 3666
rect 25342 3614 25394 3666
rect 27694 3614 27746 3666
rect 28590 3614 28642 3666
rect 29262 3614 29314 3666
rect 32174 3614 32226 3666
rect 33182 3614 33234 3666
rect 35870 3614 35922 3666
rect 37102 3614 37154 3666
rect 42030 3614 42082 3666
rect 3054 3502 3106 3554
rect 4734 3502 4786 3554
rect 5854 3502 5906 3554
rect 7870 3502 7922 3554
rect 9774 3502 9826 3554
rect 11566 3502 11618 3554
rect 13582 3502 13634 3554
rect 15598 3502 15650 3554
rect 17614 3502 17666 3554
rect 19406 3502 19458 3554
rect 27358 3502 27410 3554
rect 27582 3502 27634 3554
rect 27806 3502 27858 3554
rect 28030 3502 28082 3554
rect 31390 3502 31442 3554
rect 31838 3502 31890 3554
rect 32398 3502 32450 3554
rect 35310 3502 35362 3554
rect 39118 3502 39170 3554
rect 39566 3502 39618 3554
rect 39790 3502 39842 3554
rect 40910 3502 40962 3554
rect 41358 3502 41410 3554
rect 41582 3502 41634 3554
rect 3838 3390 3890 3442
rect 8766 3390 8818 3442
rect 22542 3390 22594 3442
rect 26350 3390 26402 3442
rect 30270 3390 30322 3442
rect 34526 3390 34578 3442
rect 38110 3390 38162 3442
rect 39342 3390 39394 3442
rect 41470 3390 41522 3442
rect 32510 3278 32562 3330
rect 35422 3278 35474 3330
rect 40126 3278 40178 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 21952 43200 22064 44000
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 18396 39060 18452 39070
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 14364 24836 14420 24846
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 3276 22484 3332 22494
rect 3276 22482 3444 22484
rect 3276 22430 3278 22482
rect 3330 22430 3444 22482
rect 3276 22428 3444 22430
rect 3276 22418 3332 22428
rect 3388 22372 3444 22428
rect 3388 22306 3444 22316
rect 8428 22372 8484 22382
rect 1932 22258 1988 22270
rect 1932 22206 1934 22258
rect 1986 22206 1988 22258
rect 1820 22036 1876 22046
rect 1932 22036 1988 22206
rect 1876 21980 1988 22036
rect 1820 21810 1876 21980
rect 1820 21758 1822 21810
rect 1874 21758 1876 21810
rect 1820 21746 1876 21758
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1596 20916 1652 20926
rect 1148 4228 1204 4238
rect 1148 800 1204 4172
rect 1596 2660 1652 20860
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1596 2594 1652 2604
rect 1708 18340 1764 18350
rect 1708 2436 1764 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 6748 15876 6804 15886
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 6412 13860 6468 13870
rect 3948 13748 4004 13758
rect 2940 13636 2996 13646
rect 2044 12628 2100 12638
rect 1932 9602 1988 9614
rect 1932 9550 1934 9602
rect 1986 9550 1988 9602
rect 1820 9492 1876 9502
rect 1820 7698 1876 9436
rect 1932 9156 1988 9550
rect 1932 9090 1988 9100
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 7634 1876 7646
rect 1932 8260 1988 8270
rect 1932 6802 1988 8204
rect 1932 6750 1934 6802
rect 1986 6750 1988 6802
rect 1932 6738 1988 6750
rect 2044 6132 2100 12572
rect 2828 11956 2884 11966
rect 2716 10836 2772 10846
rect 2716 10742 2772 10780
rect 2380 10050 2436 10062
rect 2380 9998 2382 10050
rect 2434 9998 2436 10050
rect 2380 9938 2436 9998
rect 2380 9886 2382 9938
rect 2434 9886 2436 9938
rect 2380 9874 2436 9886
rect 2828 9938 2884 11900
rect 2828 9886 2830 9938
rect 2882 9886 2884 9938
rect 2828 9874 2884 9886
rect 2604 9380 2660 9390
rect 2156 8930 2212 8942
rect 2492 8932 2548 8942
rect 2156 8878 2158 8930
rect 2210 8878 2212 8930
rect 2156 8372 2212 8878
rect 2156 8306 2212 8316
rect 2268 8930 2548 8932
rect 2268 8878 2494 8930
rect 2546 8878 2548 8930
rect 2268 8876 2548 8878
rect 2156 8036 2212 8046
rect 2156 6132 2212 7980
rect 2268 7924 2324 8876
rect 2492 8866 2548 8876
rect 2604 8428 2660 9324
rect 2268 7698 2324 7868
rect 2268 7646 2270 7698
rect 2322 7646 2324 7698
rect 2268 7634 2324 7646
rect 2380 8372 2660 8428
rect 2380 6690 2436 8372
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7252 2548 7982
rect 2828 8036 2884 8046
rect 2828 7942 2884 7980
rect 2492 7186 2548 7196
rect 2604 7812 2660 7822
rect 2380 6638 2382 6690
rect 2434 6638 2436 6690
rect 2380 6626 2436 6638
rect 2268 6132 2324 6142
rect 2156 6130 2324 6132
rect 2156 6078 2270 6130
rect 2322 6078 2324 6130
rect 2156 6076 2324 6078
rect 2044 6066 2100 6076
rect 2268 6066 2324 6076
rect 1820 5794 1876 5806
rect 1820 5742 1822 5794
rect 1874 5742 1876 5794
rect 1820 4676 1876 5742
rect 2156 5682 2212 5694
rect 2156 5630 2158 5682
rect 2210 5630 2212 5682
rect 2156 5234 2212 5630
rect 2156 5182 2158 5234
rect 2210 5182 2212 5234
rect 2156 5170 2212 5182
rect 2604 5234 2660 7756
rect 2716 7700 2772 7710
rect 2716 7606 2772 7644
rect 2716 6466 2772 6478
rect 2716 6414 2718 6466
rect 2770 6414 2772 6466
rect 2716 6244 2772 6414
rect 2716 6130 2772 6188
rect 2716 6078 2718 6130
rect 2770 6078 2772 6130
rect 2716 6066 2772 6078
rect 2940 5682 2996 13580
rect 3612 11172 3668 11182
rect 3164 10500 3220 10510
rect 3164 10498 3332 10500
rect 3164 10446 3166 10498
rect 3218 10446 3332 10498
rect 3164 10444 3332 10446
rect 3164 10434 3220 10444
rect 3164 10050 3220 10062
rect 3164 9998 3166 10050
rect 3218 9998 3220 10050
rect 3164 9828 3220 9998
rect 3276 10052 3332 10444
rect 3276 9986 3332 9996
rect 3500 10498 3556 10510
rect 3500 10446 3502 10498
rect 3554 10446 3556 10498
rect 3500 9828 3556 10446
rect 3612 10052 3668 11116
rect 3612 9986 3668 9996
rect 3164 9772 3556 9828
rect 3836 9828 3892 9838
rect 3164 9602 3220 9772
rect 3164 9550 3166 9602
rect 3218 9550 3220 9602
rect 3164 9380 3220 9550
rect 3612 9602 3668 9614
rect 3612 9550 3614 9602
rect 3666 9550 3668 9602
rect 3612 9492 3668 9550
rect 3612 9426 3668 9436
rect 3836 9604 3892 9772
rect 3164 9324 3556 9380
rect 3500 9268 3556 9324
rect 3500 9212 3668 9268
rect 3052 8932 3108 8942
rect 3052 8838 3108 8876
rect 3388 8930 3444 8942
rect 3388 8878 3390 8930
rect 3442 8878 3444 8930
rect 3388 8818 3444 8878
rect 3388 8766 3390 8818
rect 3442 8766 3444 8818
rect 3388 8754 3444 8766
rect 3500 8820 3556 8830
rect 3388 8482 3444 8494
rect 3388 8430 3390 8482
rect 3442 8430 3444 8482
rect 3164 8372 3220 8382
rect 3052 8260 3108 8270
rect 3052 7698 3108 8204
rect 3052 7646 3054 7698
rect 3106 7646 3108 7698
rect 3052 7634 3108 7646
rect 3164 6692 3220 8316
rect 3388 8370 3444 8430
rect 3388 8318 3390 8370
rect 3442 8318 3444 8370
rect 3388 8306 3444 8318
rect 3164 6626 3220 6636
rect 3276 6692 3332 6702
rect 3500 6692 3556 8764
rect 3612 7700 3668 9212
rect 3836 9266 3892 9548
rect 3836 9214 3838 9266
rect 3890 9214 3892 9266
rect 3836 9202 3892 9214
rect 3724 9156 3780 9166
rect 3724 7812 3780 9100
rect 3836 8372 3892 8382
rect 3948 8372 4004 13692
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 5964 13300 6020 13310
rect 5964 12738 6020 13244
rect 6412 13074 6468 13804
rect 6748 13634 6804 15820
rect 8428 14980 8484 22316
rect 11340 20692 11396 20702
rect 10108 15204 10164 15214
rect 8428 14914 8484 14924
rect 9660 15092 9716 15102
rect 9660 14644 9716 15036
rect 9548 14642 9716 14644
rect 9548 14590 9662 14642
rect 9714 14590 9716 14642
rect 9548 14588 9716 14590
rect 9212 14306 9268 14318
rect 9212 14254 9214 14306
rect 9266 14254 9268 14306
rect 9100 13860 9156 13870
rect 6748 13582 6750 13634
rect 6802 13582 6804 13634
rect 6748 13522 6804 13582
rect 6748 13470 6750 13522
rect 6802 13470 6804 13522
rect 6748 13458 6804 13470
rect 7196 13634 7252 13646
rect 7196 13582 7198 13634
rect 7250 13582 7252 13634
rect 7196 13300 7252 13582
rect 7644 13634 7700 13646
rect 7644 13582 7646 13634
rect 7698 13582 7700 13634
rect 7420 13522 7476 13534
rect 7420 13470 7422 13522
rect 7474 13470 7476 13522
rect 7420 13300 7476 13470
rect 7644 13522 7700 13582
rect 7644 13470 7646 13522
rect 7698 13470 7700 13522
rect 7644 13458 7700 13470
rect 8092 13634 8148 13646
rect 8092 13582 8094 13634
rect 8146 13582 8148 13634
rect 7420 13244 8036 13300
rect 7196 13234 7252 13244
rect 6412 13022 6414 13074
rect 6466 13022 6468 13074
rect 6412 13010 6468 13022
rect 7196 13074 7252 13086
rect 7196 13022 7198 13074
rect 7250 13022 7252 13074
rect 5964 12686 5966 12738
rect 6018 12686 6020 12738
rect 5964 12292 6020 12686
rect 5516 12236 6020 12292
rect 4732 12068 4788 12078
rect 4732 12066 4900 12068
rect 4732 12014 4734 12066
rect 4786 12014 4900 12066
rect 4732 12012 4900 12014
rect 4732 12002 4788 12012
rect 4284 11956 4340 11966
rect 4060 11172 4116 11182
rect 4060 11078 4116 11116
rect 4284 10836 4340 11900
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4844 11788 4900 12012
rect 5068 12066 5124 12078
rect 5068 12014 5070 12066
rect 5122 12014 5124 12066
rect 4844 11732 5012 11788
rect 4476 11722 4740 11732
rect 4508 11172 4564 11182
rect 4508 11078 4564 11116
rect 4956 11170 5012 11732
rect 4956 11118 4958 11170
rect 5010 11118 5012 11170
rect 4956 11060 5012 11118
rect 4956 10994 5012 11004
rect 4396 10836 4452 10846
rect 4284 10834 4452 10836
rect 4284 10782 4398 10834
rect 4450 10782 4452 10834
rect 4284 10780 4452 10782
rect 5068 10836 5124 12014
rect 5292 11172 5348 11182
rect 5180 10836 5236 10846
rect 5068 10780 5180 10836
rect 4396 10770 4452 10780
rect 4060 10500 4116 10510
rect 4060 10406 4116 10444
rect 4844 10498 4900 10510
rect 4844 10446 4846 10498
rect 4898 10446 4900 10498
rect 4284 10388 4340 10398
rect 4172 9604 4228 9614
rect 4172 9510 4228 9548
rect 4284 9156 4340 10332
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4508 10052 4564 10062
rect 4508 9938 4564 9996
rect 4508 9886 4510 9938
rect 4562 9886 4564 9938
rect 4172 9100 4340 9156
rect 4396 9380 4452 9390
rect 4060 8932 4116 8942
rect 4060 8482 4116 8876
rect 4172 8708 4228 9100
rect 4284 8932 4340 8942
rect 4396 8932 4452 9324
rect 4340 8876 4452 8932
rect 4284 8800 4340 8876
rect 4508 8818 4564 9886
rect 4844 9716 4900 10446
rect 5068 9940 5124 9950
rect 5068 9846 5124 9884
rect 4844 9156 4900 9660
rect 4844 9090 4900 9100
rect 4732 8932 4788 8942
rect 4732 8930 4900 8932
rect 4732 8878 4734 8930
rect 4786 8878 4900 8930
rect 4732 8876 4900 8878
rect 4732 8866 4788 8876
rect 4508 8766 4510 8818
rect 4562 8766 4564 8818
rect 4508 8754 4564 8766
rect 4172 8652 4340 8708
rect 4060 8430 4062 8482
rect 4114 8430 4116 8482
rect 4060 8418 4116 8430
rect 3836 8370 4004 8372
rect 3836 8318 3838 8370
rect 3890 8318 4004 8370
rect 3836 8316 4004 8318
rect 3836 8306 3892 8316
rect 4172 8260 4228 8270
rect 4172 8166 4228 8204
rect 3724 7756 3892 7812
rect 3612 7634 3668 7644
rect 3724 7588 3780 7598
rect 3724 7494 3780 7532
rect 3612 7362 3668 7374
rect 3612 7310 3614 7362
rect 3666 7310 3668 7362
rect 3612 6804 3668 7310
rect 3612 6738 3668 6748
rect 3276 6690 3556 6692
rect 3276 6638 3278 6690
rect 3330 6638 3556 6690
rect 3276 6636 3556 6638
rect 3276 6626 3332 6636
rect 3724 6466 3780 6478
rect 3724 6414 3726 6466
rect 3778 6414 3780 6466
rect 3164 6132 3220 6142
rect 3164 6038 3220 6076
rect 3612 5796 3668 5806
rect 2940 5630 2942 5682
rect 2994 5630 2996 5682
rect 2940 5618 2996 5630
rect 3500 5794 3668 5796
rect 3500 5742 3614 5794
rect 3666 5742 3668 5794
rect 3500 5740 3668 5742
rect 3164 5348 3220 5358
rect 2604 5182 2606 5234
rect 2658 5182 2660 5234
rect 2604 5170 2660 5182
rect 2940 5236 2996 5246
rect 1820 4610 1876 4620
rect 2940 4338 2996 5180
rect 3164 5234 3220 5292
rect 3164 5182 3166 5234
rect 3218 5182 3220 5234
rect 3164 5170 3220 5182
rect 2940 4286 2942 4338
rect 2994 4286 2996 4338
rect 2940 4274 2996 4286
rect 3052 4898 3108 4910
rect 3052 4846 3054 4898
rect 3106 4846 3108 4898
rect 1932 4228 1988 4238
rect 1932 4134 1988 4172
rect 1708 2370 1764 2380
rect 2492 3666 2548 3678
rect 2492 3614 2494 3666
rect 2546 3614 2548 3666
rect 2492 800 2548 3614
rect 3052 3554 3108 4846
rect 3052 3502 3054 3554
rect 3106 3502 3108 3554
rect 3052 3490 3108 3502
rect 3500 2996 3556 5740
rect 3612 5730 3668 5740
rect 3612 5124 3668 5134
rect 3612 4450 3668 5068
rect 3612 4398 3614 4450
rect 3666 4398 3668 4450
rect 3612 4386 3668 4398
rect 3724 4340 3780 6414
rect 3836 5460 3892 7756
rect 4284 7586 4340 8652
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4732 8372 4788 8382
rect 4732 8258 4788 8316
rect 4732 8206 4734 8258
rect 4786 8206 4788 8258
rect 4284 7534 4286 7586
rect 4338 7534 4340 7586
rect 4284 7522 4340 7534
rect 4508 7812 4564 7822
rect 4396 7476 4452 7486
rect 4396 7382 4452 7420
rect 4508 7252 4564 7756
rect 4732 7812 4788 8206
rect 4844 8260 4900 8876
rect 5068 8596 5124 8606
rect 4844 8194 4900 8204
rect 4956 8484 5012 8494
rect 4844 8036 4900 8046
rect 4956 8036 5012 8428
rect 5068 8372 5124 8540
rect 5068 8306 5124 8316
rect 5180 8260 5236 10780
rect 5292 10498 5348 11116
rect 5292 10446 5294 10498
rect 5346 10446 5348 10498
rect 5292 9268 5348 10446
rect 5292 9202 5348 9212
rect 5404 9156 5460 9166
rect 5404 9062 5460 9100
rect 5292 8818 5348 8830
rect 5292 8766 5294 8818
rect 5346 8766 5348 8818
rect 5292 8484 5348 8766
rect 5292 8418 5348 8428
rect 5180 8204 5460 8260
rect 4844 8034 5012 8036
rect 4844 7982 4846 8034
rect 4898 7982 5012 8034
rect 4844 7980 5012 7982
rect 5068 8034 5124 8046
rect 5068 7982 5070 8034
rect 5122 7982 5124 8034
rect 4844 7970 4900 7980
rect 5068 7812 5124 7982
rect 4732 7756 5012 7812
rect 4620 7700 4676 7710
rect 4732 7700 4788 7756
rect 4676 7644 4788 7700
rect 4620 7634 4676 7644
rect 4956 7586 5012 7756
rect 5068 7746 5124 7756
rect 5180 8036 5236 8046
rect 4956 7534 4958 7586
rect 5010 7534 5012 7586
rect 4956 7522 5012 7534
rect 5068 7588 5124 7598
rect 5180 7588 5236 7980
rect 5068 7586 5236 7588
rect 5068 7534 5070 7586
rect 5122 7534 5236 7586
rect 5068 7532 5236 7534
rect 5068 7522 5124 7532
rect 5292 7474 5348 7486
rect 5292 7422 5294 7474
rect 5346 7422 5348 7474
rect 5180 7364 5236 7374
rect 4508 7196 4900 7252
rect 4844 7140 4900 7196
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4844 7074 4900 7084
rect 4476 7018 4740 7028
rect 4172 6578 4228 6590
rect 4172 6526 4174 6578
rect 4226 6526 4228 6578
rect 4172 6468 4228 6526
rect 4844 6580 4900 6590
rect 4844 6486 4900 6524
rect 4172 6402 4228 6412
rect 4284 6466 4340 6478
rect 4284 6414 4286 6466
rect 4338 6414 4340 6466
rect 3836 5394 3892 5404
rect 3948 5908 4004 5918
rect 3948 5348 4004 5852
rect 4060 5796 4116 5806
rect 4060 5794 4228 5796
rect 4060 5742 4062 5794
rect 4114 5742 4228 5794
rect 4060 5740 4228 5742
rect 4060 5730 4116 5740
rect 3948 5216 4004 5292
rect 4060 5572 4116 5582
rect 4060 5122 4116 5516
rect 4060 5070 4062 5122
rect 4114 5070 4116 5122
rect 3948 4900 4004 4910
rect 3724 4274 3780 4284
rect 3836 4898 4004 4900
rect 3836 4846 3950 4898
rect 4002 4846 4004 4898
rect 3836 4844 4004 4846
rect 3836 4116 3892 4844
rect 3948 4834 4004 4844
rect 4060 4788 4116 5070
rect 4060 4722 4116 4732
rect 3948 4452 4004 4462
rect 3948 4358 4004 4396
rect 3836 4050 3892 4060
rect 3500 2930 3556 2940
rect 3836 3442 3892 3454
rect 3836 3390 3838 3442
rect 3890 3390 3892 3442
rect 3836 800 3892 3390
rect 4172 3332 4228 5740
rect 4284 3556 4340 6414
rect 4956 6466 5012 6478
rect 4956 6414 4958 6466
rect 5010 6414 5012 6466
rect 4620 6244 4676 6254
rect 4620 6130 4676 6188
rect 4620 6078 4622 6130
rect 4674 6078 4676 6130
rect 4620 6066 4676 6078
rect 4956 6132 5012 6414
rect 4956 6066 5012 6076
rect 4732 5908 4788 5918
rect 4732 5906 5012 5908
rect 4732 5854 4734 5906
rect 4786 5854 5012 5906
rect 4732 5852 5012 5854
rect 4732 5842 4788 5852
rect 4844 5684 4900 5694
rect 4844 5590 4900 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4508 5348 4564 5358
rect 4508 4450 4564 5292
rect 4956 5124 5012 5852
rect 5180 5796 5236 7308
rect 5292 7028 5348 7422
rect 5292 6962 5348 6972
rect 5180 5730 5236 5740
rect 5292 6692 5348 6702
rect 5292 5572 5348 6636
rect 5404 6244 5460 8204
rect 5516 6692 5572 12236
rect 6076 12180 6132 12190
rect 5964 12178 6132 12180
rect 5964 12126 6078 12178
rect 6130 12126 6132 12178
rect 5964 12124 6132 12126
rect 5628 12068 5684 12078
rect 5628 12066 5908 12068
rect 5628 12014 5630 12066
rect 5682 12014 5908 12066
rect 5628 12012 5908 12014
rect 5628 12002 5684 12012
rect 5852 11956 5908 12012
rect 5740 10500 5796 10510
rect 5740 10406 5796 10444
rect 5628 10052 5684 10062
rect 5628 9602 5684 9996
rect 5628 9550 5630 9602
rect 5682 9550 5684 9602
rect 5628 8372 5684 9550
rect 5628 8306 5684 8316
rect 5740 9380 5796 9390
rect 5628 8148 5684 8186
rect 5628 8082 5684 8092
rect 5740 7700 5796 9324
rect 5852 8260 5908 11900
rect 5964 9940 6020 12124
rect 6076 12114 6132 12124
rect 6300 12180 6356 12190
rect 6076 11284 6132 11294
rect 6076 11190 6132 11228
rect 6188 11172 6244 11182
rect 6188 11078 6244 11116
rect 6300 10948 6356 12124
rect 6860 12066 6916 12078
rect 6860 12014 6862 12066
rect 6914 12014 6916 12066
rect 6860 11506 6916 12014
rect 7196 11844 7252 13022
rect 7196 11778 7252 11788
rect 6860 11454 6862 11506
rect 6914 11454 6916 11506
rect 6860 11442 6916 11454
rect 7084 11396 7140 11406
rect 7756 11396 7812 11406
rect 7084 11394 7812 11396
rect 7084 11342 7086 11394
rect 7138 11342 7758 11394
rect 7810 11342 7812 11394
rect 7084 11340 7812 11342
rect 7084 11330 7140 11340
rect 7756 11330 7812 11340
rect 6748 11282 6804 11294
rect 6748 11230 6750 11282
rect 6802 11230 6804 11282
rect 6748 11172 6804 11230
rect 6748 11106 6804 11116
rect 7644 11170 7700 11182
rect 7644 11118 7646 11170
rect 7698 11118 7700 11170
rect 5964 9874 6020 9884
rect 6188 10892 6356 10948
rect 6972 11060 7028 11070
rect 6076 9716 6132 9726
rect 6076 9622 6132 9660
rect 6188 9380 6244 10892
rect 6300 10724 6356 10734
rect 6300 10630 6356 10668
rect 6860 10612 6916 10622
rect 6636 10556 6860 10612
rect 6636 9938 6692 10556
rect 6860 10518 6916 10556
rect 6748 10386 6804 10398
rect 6748 10334 6750 10386
rect 6802 10334 6804 10386
rect 6748 10052 6804 10334
rect 6748 9986 6804 9996
rect 6636 9886 6638 9938
rect 6690 9886 6692 9938
rect 6636 9874 6692 9886
rect 6972 9828 7028 11004
rect 7644 11060 7700 11118
rect 7644 10994 7700 11004
rect 7868 11170 7924 11182
rect 7868 11118 7870 11170
rect 7922 11118 7924 11170
rect 7868 11060 7924 11118
rect 7644 10724 7700 10734
rect 7420 10722 7700 10724
rect 7420 10670 7646 10722
rect 7698 10670 7700 10722
rect 7420 10668 7700 10670
rect 7420 10612 7476 10668
rect 7644 10658 7700 10668
rect 5964 9324 6244 9380
rect 6748 9772 7028 9828
rect 7308 10556 7476 10612
rect 5964 9154 6020 9324
rect 5964 9102 5966 9154
rect 6018 9102 6020 9154
rect 5964 8596 6020 9102
rect 6076 9156 6132 9166
rect 6132 9100 6244 9156
rect 6076 9024 6132 9100
rect 5964 8530 6020 8540
rect 6188 8484 6244 9100
rect 6300 9044 6356 9054
rect 6300 8950 6356 8988
rect 6748 9042 6804 9772
rect 7196 9492 7252 9502
rect 6748 8990 6750 9042
rect 6802 8990 6804 9042
rect 6524 8484 6580 8494
rect 6188 8482 6580 8484
rect 6188 8430 6526 8482
rect 6578 8430 6580 8482
rect 6188 8428 6580 8430
rect 6524 8418 6580 8428
rect 5964 8260 6020 8270
rect 6748 8260 6804 8990
rect 6860 9154 6916 9166
rect 6860 9102 6862 9154
rect 6914 9102 6916 9154
rect 6860 8932 6916 9102
rect 7084 9156 7140 9166
rect 7084 9062 7140 9100
rect 6860 8866 6916 8876
rect 5852 8258 6020 8260
rect 5852 8206 5966 8258
rect 6018 8206 6020 8258
rect 5852 8204 6020 8206
rect 5964 8194 6020 8204
rect 6524 8204 6804 8260
rect 5852 8036 5908 8046
rect 5852 7942 5908 7980
rect 5740 7644 5908 7700
rect 5852 7586 5908 7644
rect 5852 7534 5854 7586
rect 5906 7534 5908 7586
rect 5852 7522 5908 7534
rect 5740 7474 5796 7486
rect 5740 7422 5742 7474
rect 5794 7422 5796 7474
rect 5740 7140 5796 7422
rect 5852 7252 5908 7262
rect 5852 7158 5908 7196
rect 5740 7074 5796 7084
rect 6076 7140 6132 7150
rect 5516 6636 5796 6692
rect 5628 6468 5684 6478
rect 5628 6374 5684 6412
rect 5404 6188 5684 6244
rect 5516 6020 5572 6030
rect 5516 5926 5572 5964
rect 5628 5796 5684 6188
rect 5740 6020 5796 6636
rect 5964 6580 6020 6590
rect 5964 6486 6020 6524
rect 5852 6466 5908 6478
rect 5852 6414 5854 6466
rect 5906 6414 5908 6466
rect 5852 6356 5908 6414
rect 5852 6300 6020 6356
rect 5740 5926 5796 5964
rect 5964 5796 6020 6300
rect 5628 5740 6020 5796
rect 5292 5506 5348 5516
rect 5404 5682 5460 5694
rect 5404 5630 5406 5682
rect 5458 5630 5460 5682
rect 5404 5236 5460 5630
rect 5404 5170 5460 5180
rect 5740 5124 5796 5134
rect 4956 5068 5124 5124
rect 4620 5012 4676 5022
rect 5068 5012 5124 5068
rect 5740 5030 5796 5068
rect 5068 4956 5348 5012
rect 4620 4918 4676 4956
rect 4956 4900 5012 4910
rect 4956 4806 5012 4844
rect 4732 4564 4788 4574
rect 4732 4470 4788 4508
rect 4508 4398 4510 4450
rect 4562 4398 4564 4450
rect 4508 4386 4564 4398
rect 5292 4340 5348 4956
rect 5852 4452 5908 4462
rect 5404 4340 5460 4350
rect 5292 4338 5460 4340
rect 5292 4286 5406 4338
rect 5458 4286 5460 4338
rect 5292 4284 5460 4286
rect 5404 4274 5460 4284
rect 5180 4228 5236 4238
rect 4844 4114 4900 4126
rect 4844 4062 4846 4114
rect 4898 4062 4900 4114
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4732 3556 4788 3566
rect 4284 3554 4788 3556
rect 4284 3502 4734 3554
rect 4786 3502 4788 3554
rect 4284 3500 4788 3502
rect 4732 3490 4788 3500
rect 4844 3556 4900 4062
rect 4844 3490 4900 3500
rect 4172 3266 4228 3276
rect 5180 800 5236 4172
rect 5852 3554 5908 4396
rect 5964 4116 6020 5740
rect 6076 5346 6132 7084
rect 6524 7140 6580 8204
rect 6860 8148 6916 8158
rect 7196 8148 7252 9436
rect 7308 9044 7364 10556
rect 7532 10500 7588 10510
rect 7868 10500 7924 11004
rect 7532 10498 7924 10500
rect 7532 10446 7534 10498
rect 7586 10446 7924 10498
rect 7532 10444 7924 10446
rect 7308 8978 7364 8988
rect 7420 10386 7476 10398
rect 7420 10334 7422 10386
rect 7474 10334 7476 10386
rect 7420 10052 7476 10334
rect 7420 8820 7476 9996
rect 7532 9154 7588 10444
rect 7980 10388 8036 13244
rect 8092 11396 8148 13582
rect 8652 13634 8708 13646
rect 8652 13582 8654 13634
rect 8706 13582 8708 13634
rect 8540 12740 8596 12750
rect 8092 11282 8148 11340
rect 8092 11230 8094 11282
rect 8146 11230 8148 11282
rect 8092 11218 8148 11230
rect 8204 11844 8260 11854
rect 8204 10948 8260 11788
rect 7868 10332 8036 10388
rect 8092 10892 8260 10948
rect 8428 11396 8484 11406
rect 7532 9102 7534 9154
rect 7586 9102 7588 9154
rect 7532 9090 7588 9102
rect 7644 9604 7700 9614
rect 7420 8708 7476 8764
rect 6860 8146 7028 8148
rect 6860 8094 6862 8146
rect 6914 8094 7028 8146
rect 6860 8092 7028 8094
rect 6860 8082 6916 8092
rect 6636 8036 6692 8046
rect 6636 7942 6692 7980
rect 6748 7812 6804 7822
rect 6748 7698 6804 7756
rect 6748 7646 6750 7698
rect 6802 7646 6804 7698
rect 6748 7634 6804 7646
rect 6972 7588 7028 8092
rect 7196 8082 7252 8092
rect 7308 8652 7476 8708
rect 6972 7494 7028 7532
rect 7084 8036 7140 8046
rect 6524 7074 6580 7084
rect 6636 7474 6692 7486
rect 6636 7422 6638 7474
rect 6690 7422 6692 7474
rect 6300 7028 6356 7038
rect 6300 5906 6356 6972
rect 6524 6804 6580 6814
rect 6524 6710 6580 6748
rect 6636 6468 6692 7422
rect 7084 7474 7140 7980
rect 7084 7422 7086 7474
rect 7138 7422 7140 7474
rect 7084 7410 7140 7422
rect 6860 7364 6916 7374
rect 6860 7270 6916 7308
rect 6636 6402 6692 6412
rect 6748 6132 6804 6142
rect 6748 6038 6804 6076
rect 6972 6020 7028 6030
rect 6972 5926 7028 5964
rect 6300 5854 6302 5906
rect 6354 5854 6356 5906
rect 6300 5842 6356 5854
rect 6524 5908 6580 5918
rect 6524 5814 6580 5852
rect 6636 5794 6692 5806
rect 6636 5742 6638 5794
rect 6690 5742 6692 5794
rect 6076 5294 6078 5346
rect 6130 5294 6132 5346
rect 6076 5282 6132 5294
rect 6300 5572 6356 5582
rect 6300 5234 6356 5516
rect 6300 5182 6302 5234
rect 6354 5182 6356 5234
rect 6300 5170 6356 5182
rect 6636 5236 6692 5742
rect 7308 5684 7364 8652
rect 7644 8596 7700 9548
rect 7756 9044 7812 9054
rect 7868 9044 7924 10332
rect 7980 9268 8036 9278
rect 7980 9174 8036 9212
rect 7868 8988 8036 9044
rect 7756 8950 7812 8988
rect 7756 8596 7812 8606
rect 7644 8540 7756 8596
rect 7756 8258 7812 8540
rect 7756 8206 7758 8258
rect 7810 8206 7812 8258
rect 7756 8194 7812 8206
rect 7420 8146 7476 8158
rect 7420 8094 7422 8146
rect 7474 8094 7476 8146
rect 7420 7700 7476 8094
rect 7868 8148 7924 8158
rect 7532 8036 7588 8046
rect 7532 7942 7588 7980
rect 7420 7634 7476 7644
rect 7868 7698 7924 8092
rect 7868 7646 7870 7698
rect 7922 7646 7924 7698
rect 7868 7634 7924 7646
rect 7756 7362 7812 7374
rect 7756 7310 7758 7362
rect 7810 7310 7812 7362
rect 7756 6692 7812 7310
rect 7756 6626 7812 6636
rect 7756 5684 7812 5694
rect 7308 5618 7364 5628
rect 7644 5682 7812 5684
rect 7644 5630 7758 5682
rect 7810 5630 7812 5682
rect 7644 5628 7812 5630
rect 6636 5170 6692 5180
rect 6860 5234 6916 5246
rect 6860 5182 6862 5234
rect 6914 5182 6916 5234
rect 6860 4788 6916 5182
rect 7644 5012 7700 5628
rect 7756 5618 7812 5628
rect 7868 5684 7924 5694
rect 7644 4946 7700 4956
rect 6860 4722 6916 4732
rect 7756 4900 7812 4910
rect 7756 4338 7812 4844
rect 7756 4286 7758 4338
rect 7810 4286 7812 4338
rect 7756 4274 7812 4286
rect 6076 4228 6132 4238
rect 6076 4134 6132 4172
rect 7308 4228 7364 4238
rect 7308 4134 7364 4172
rect 5964 4050 6020 4060
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5852 3490 5908 3502
rect 6524 3666 6580 3678
rect 6524 3614 6526 3666
rect 6578 3614 6580 3666
rect 6524 800 6580 3614
rect 7868 3554 7924 5628
rect 7980 5572 8036 8988
rect 8092 8932 8148 10892
rect 8428 10834 8484 11340
rect 8428 10782 8430 10834
rect 8482 10782 8484 10834
rect 8428 10770 8484 10782
rect 8316 10612 8372 10622
rect 8316 10518 8372 10556
rect 8428 10388 8484 10398
rect 8204 10386 8484 10388
rect 8204 10334 8430 10386
rect 8482 10334 8484 10386
rect 8204 10332 8484 10334
rect 8204 9042 8260 10332
rect 8428 10322 8484 10332
rect 8204 8990 8206 9042
rect 8258 8990 8260 9042
rect 8204 8978 8260 8990
rect 8540 9044 8596 12684
rect 8652 11844 8708 13582
rect 8988 13636 9044 13646
rect 8988 13542 9044 13580
rect 8876 13522 8932 13534
rect 8876 13470 8878 13522
rect 8930 13470 8932 13522
rect 8876 12068 8932 13470
rect 8988 12068 9044 12078
rect 8876 12066 9044 12068
rect 8876 12014 8990 12066
rect 9042 12014 9044 12066
rect 8876 12012 9044 12014
rect 8652 11778 8708 11788
rect 8652 11284 8708 11294
rect 8652 11190 8708 11228
rect 8988 11282 9044 12012
rect 8988 11230 8990 11282
rect 9042 11230 9044 11282
rect 8876 11170 8932 11182
rect 8876 11118 8878 11170
rect 8930 11118 8932 11170
rect 8876 11060 8932 11118
rect 8876 10994 8932 11004
rect 8988 10948 9044 11230
rect 8988 10882 9044 10892
rect 8988 10498 9044 10510
rect 8988 10446 8990 10498
rect 9042 10446 9044 10498
rect 8988 9940 9044 10446
rect 8988 9874 9044 9884
rect 8764 9714 8820 9726
rect 8764 9662 8766 9714
rect 8818 9662 8820 9714
rect 8764 9268 8820 9662
rect 8764 9202 8820 9212
rect 9100 9268 9156 13804
rect 9212 13522 9268 14254
rect 9212 13470 9214 13522
rect 9266 13470 9268 13522
rect 9212 13458 9268 13470
rect 9324 12850 9380 12862
rect 9324 12798 9326 12850
rect 9378 12798 9380 12850
rect 9324 12292 9380 12798
rect 9324 12226 9380 12236
rect 9436 12404 9492 12414
rect 9436 11844 9492 12348
rect 9324 11788 9492 11844
rect 9100 9202 9156 9212
rect 9212 9716 9268 9726
rect 8876 9156 8932 9166
rect 8876 9062 8932 9100
rect 8540 8988 8820 9044
rect 8092 5906 8148 8876
rect 8204 8372 8260 8382
rect 8204 8258 8260 8316
rect 8540 8370 8596 8988
rect 8652 8820 8708 8830
rect 8652 8726 8708 8764
rect 8540 8318 8542 8370
rect 8594 8318 8596 8370
rect 8540 8306 8596 8318
rect 8652 8484 8708 8494
rect 8204 8206 8206 8258
rect 8258 8206 8260 8258
rect 8204 8194 8260 8206
rect 8092 5854 8094 5906
rect 8146 5854 8148 5906
rect 8092 5842 8148 5854
rect 8428 8034 8484 8046
rect 8428 7982 8430 8034
rect 8482 7982 8484 8034
rect 7980 5506 8036 5516
rect 8316 5794 8372 5806
rect 8316 5742 8318 5794
rect 8370 5742 8372 5794
rect 8316 5572 8372 5742
rect 8428 5684 8484 7982
rect 8652 7924 8708 8428
rect 8764 8258 8820 8988
rect 8988 8932 9044 8942
rect 8988 8838 9044 8876
rect 8764 8206 8766 8258
rect 8818 8206 8820 8258
rect 8764 8194 8820 8206
rect 8876 8820 8932 8830
rect 8876 8036 8932 8764
rect 9212 8820 9268 9660
rect 9212 8754 9268 8764
rect 8540 7868 8708 7924
rect 8764 7980 8932 8036
rect 8988 8258 9044 8270
rect 8988 8206 8990 8258
rect 9042 8206 9044 8258
rect 8540 7474 8596 7868
rect 8540 7422 8542 7474
rect 8594 7422 8596 7474
rect 8540 7410 8596 7422
rect 8764 7474 8820 7980
rect 8876 7698 8932 7710
rect 8876 7646 8878 7698
rect 8930 7646 8932 7698
rect 8876 7588 8932 7646
rect 8876 7522 8932 7532
rect 8764 7422 8766 7474
rect 8818 7422 8820 7474
rect 8764 7410 8820 7422
rect 8988 7474 9044 8206
rect 9100 8146 9156 8158
rect 9100 8094 9102 8146
rect 9154 8094 9156 8146
rect 9100 7924 9156 8094
rect 9100 7858 9156 7868
rect 9212 8034 9268 8046
rect 9212 7982 9214 8034
rect 9266 7982 9268 8034
rect 8988 7422 8990 7474
rect 9042 7422 9044 7474
rect 8988 7410 9044 7422
rect 8652 7364 8708 7374
rect 8652 6690 8708 7308
rect 8652 6638 8654 6690
rect 8706 6638 8708 6690
rect 8652 6626 8708 6638
rect 8876 6468 8932 6478
rect 8876 6018 8932 6412
rect 8876 5966 8878 6018
rect 8930 5966 8932 6018
rect 8876 5954 8932 5966
rect 8428 5618 8484 5628
rect 8988 5684 9044 5694
rect 8988 5682 9156 5684
rect 8988 5630 8990 5682
rect 9042 5630 9156 5682
rect 8988 5628 9156 5630
rect 8988 5618 9044 5628
rect 8316 5506 8372 5516
rect 8988 5236 9044 5246
rect 8988 5142 9044 5180
rect 9100 4564 9156 5628
rect 9212 4676 9268 7982
rect 9324 6580 9380 11788
rect 9436 9940 9492 9950
rect 9436 9826 9492 9884
rect 9436 9774 9438 9826
rect 9490 9774 9492 9826
rect 9436 9762 9492 9774
rect 9436 8372 9492 8382
rect 9436 8258 9492 8316
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 9436 8194 9492 8206
rect 9436 6804 9492 6814
rect 9436 6690 9492 6748
rect 9436 6638 9438 6690
rect 9490 6638 9492 6690
rect 9436 6626 9492 6638
rect 9324 6514 9380 6524
rect 9548 6468 9604 14588
rect 9660 14578 9716 14588
rect 10108 14642 10164 15148
rect 10108 14590 10110 14642
rect 10162 14590 10164 14642
rect 10108 14578 10164 14590
rect 11228 14754 11284 14766
rect 11228 14702 11230 14754
rect 11282 14702 11284 14754
rect 11116 14306 11172 14318
rect 11116 14254 11118 14306
rect 11170 14254 11172 14306
rect 11116 13860 11172 14254
rect 11116 13794 11172 13804
rect 9884 13634 9940 13646
rect 9884 13582 9886 13634
rect 9938 13582 9940 13634
rect 9884 12516 9940 13582
rect 10332 13636 10388 13646
rect 9884 12450 9940 12460
rect 10108 12964 10164 12974
rect 10332 12964 10388 13580
rect 10108 12962 10388 12964
rect 10108 12910 10110 12962
rect 10162 12910 10388 12962
rect 10108 12908 10388 12910
rect 11116 13636 11172 13646
rect 11228 13636 11284 14702
rect 11116 13634 11284 13636
rect 11116 13582 11118 13634
rect 11170 13582 11284 13634
rect 11116 13580 11284 13582
rect 9884 12292 9940 12302
rect 9884 12198 9940 12236
rect 9772 12068 9828 12078
rect 9660 11844 9716 11854
rect 9660 11618 9716 11788
rect 9660 11566 9662 11618
rect 9714 11566 9716 11618
rect 9660 11554 9716 11566
rect 9772 11060 9828 12012
rect 9996 11956 10052 11966
rect 9884 11954 10052 11956
rect 9884 11902 9998 11954
rect 10050 11902 10052 11954
rect 9884 11900 10052 11902
rect 9884 11506 9940 11900
rect 9996 11890 10052 11900
rect 10108 11732 10164 12908
rect 10780 12852 10836 12862
rect 10780 12850 10948 12852
rect 10780 12798 10782 12850
rect 10834 12798 10948 12850
rect 10780 12796 10948 12798
rect 10780 12786 10836 12796
rect 10668 12740 10724 12750
rect 10668 12646 10724 12684
rect 10220 12404 10276 12414
rect 10220 12178 10276 12348
rect 10556 12180 10612 12190
rect 10220 12126 10222 12178
rect 10274 12126 10276 12178
rect 10220 12114 10276 12126
rect 10444 12124 10556 12180
rect 9884 11454 9886 11506
rect 9938 11454 9940 11506
rect 9884 11442 9940 11454
rect 9996 11676 10164 11732
rect 10332 11954 10388 11966
rect 10332 11902 10334 11954
rect 10386 11902 10388 11954
rect 9884 11172 9940 11182
rect 9884 11078 9940 11116
rect 9660 11004 9828 11060
rect 9660 8484 9716 11004
rect 9996 10948 10052 11676
rect 9772 10892 10052 10948
rect 10108 11508 10164 11518
rect 9772 9940 9828 10892
rect 9884 10724 9940 10734
rect 9884 10630 9940 10668
rect 9996 10724 10052 10734
rect 10108 10724 10164 11452
rect 9996 10722 10164 10724
rect 9996 10670 9998 10722
rect 10050 10670 10164 10722
rect 9996 10668 10164 10670
rect 10332 11172 10388 11902
rect 9996 10500 10052 10668
rect 9884 10388 9940 10398
rect 9884 10294 9940 10332
rect 9772 9874 9828 9884
rect 9884 9268 9940 9278
rect 9884 9174 9940 9212
rect 9772 8818 9828 8830
rect 9772 8766 9774 8818
rect 9826 8766 9828 8818
rect 9772 8708 9828 8766
rect 9996 8708 10052 10444
rect 10332 9938 10388 11116
rect 10444 10050 10500 12124
rect 10556 12114 10612 12124
rect 10892 11788 10948 12796
rect 11116 12404 11172 13580
rect 11116 12338 11172 12348
rect 11228 12852 11284 12862
rect 11004 12180 11060 12218
rect 11004 12114 11060 12124
rect 10444 9998 10446 10050
rect 10498 9998 10500 10050
rect 10444 9986 10500 9998
rect 10556 11732 10612 11742
rect 10332 9886 10334 9938
rect 10386 9886 10388 9938
rect 10332 9874 10388 9886
rect 10108 9828 10164 9838
rect 10108 9156 10164 9772
rect 10108 9062 10164 9100
rect 10220 9602 10276 9614
rect 10220 9550 10222 9602
rect 10274 9550 10276 9602
rect 10220 9044 10276 9550
rect 10220 8978 10276 8988
rect 9772 8642 9828 8652
rect 9884 8652 10052 8708
rect 10556 8932 10612 11676
rect 10668 11732 10948 11788
rect 11116 12066 11172 12078
rect 11116 12014 11118 12066
rect 11170 12014 11172 12066
rect 11116 11844 11172 12014
rect 11116 11778 11172 11788
rect 10668 11508 10724 11732
rect 11004 11620 11060 11630
rect 11228 11620 11284 12796
rect 11004 11618 11284 11620
rect 11004 11566 11006 11618
rect 11058 11566 11284 11618
rect 11004 11564 11284 11566
rect 11004 11554 11060 11564
rect 10668 11452 10948 11508
rect 10892 11394 10948 11452
rect 10892 11342 10894 11394
rect 10946 11342 10948 11394
rect 10892 11284 10948 11342
rect 10892 10498 10948 11228
rect 11004 11172 11060 11182
rect 11004 11078 11060 11116
rect 10892 10446 10894 10498
rect 10946 10446 10948 10498
rect 10892 10434 10948 10446
rect 11116 9826 11172 11564
rect 11340 9828 11396 20636
rect 14364 16210 14420 24780
rect 18172 18564 18228 18574
rect 17276 17220 17332 17230
rect 15260 16884 15316 16894
rect 15260 16790 15316 16828
rect 14364 16158 14366 16210
rect 14418 16158 14420 16210
rect 13356 15540 13412 15550
rect 13356 15446 13412 15484
rect 14364 15540 14420 16158
rect 15372 16322 15428 16334
rect 15372 16270 15374 16322
rect 15426 16270 15428 16322
rect 14924 15876 14980 15886
rect 14924 15874 15092 15876
rect 14924 15822 14926 15874
rect 14978 15822 15092 15874
rect 14924 15820 15092 15822
rect 14924 15810 14980 15820
rect 14588 15540 14644 15550
rect 14420 15538 14644 15540
rect 14420 15486 14590 15538
rect 14642 15486 14644 15538
rect 14420 15484 14644 15486
rect 11676 15202 11732 15214
rect 11676 15150 11678 15202
rect 11730 15150 11732 15202
rect 11676 14754 11732 15150
rect 12572 15204 12628 15214
rect 12572 15110 12628 15148
rect 13020 15202 13076 15214
rect 13020 15150 13022 15202
rect 13074 15150 13076 15202
rect 13020 15148 13076 15150
rect 13916 15204 13972 15214
rect 13020 15092 13188 15148
rect 13916 15110 13972 15148
rect 14364 15148 14420 15484
rect 14588 15474 14644 15484
rect 14364 15092 14868 15148
rect 11676 14702 11678 14754
rect 11730 14702 11732 14754
rect 11676 14690 11732 14702
rect 11564 14306 11620 14318
rect 11564 14254 11566 14306
rect 11618 14254 11620 14306
rect 11564 12852 11620 14254
rect 11900 14306 11956 14318
rect 11900 14254 11902 14306
rect 11954 14254 11956 14306
rect 11676 13634 11732 13646
rect 11676 13582 11678 13634
rect 11730 13582 11732 13634
rect 11676 13076 11732 13582
rect 11900 13636 11956 14254
rect 12460 14306 12516 14318
rect 12460 14254 12462 14306
rect 12514 14254 12516 14306
rect 12012 13636 12068 13646
rect 11900 13580 12012 13636
rect 12012 13188 12068 13580
rect 12012 13132 12404 13188
rect 11676 13020 12180 13076
rect 12124 12964 12180 13020
rect 12124 12962 12292 12964
rect 12124 12910 12126 12962
rect 12178 12910 12292 12962
rect 12124 12908 12292 12910
rect 12124 12898 12180 12908
rect 12012 12852 12068 12862
rect 11564 12796 11732 12852
rect 11452 12740 11508 12750
rect 11452 11844 11508 12684
rect 11452 11778 11508 11788
rect 11564 12516 11620 12526
rect 11564 10052 11620 12460
rect 11676 11620 11732 12796
rect 12012 12758 12068 12796
rect 12236 12404 12292 12908
rect 12348 12628 12404 13132
rect 12348 12562 12404 12572
rect 12460 12516 12516 14254
rect 12908 14308 12964 14318
rect 12908 14306 13076 14308
rect 12908 14254 12910 14306
rect 12962 14254 13076 14306
rect 12908 14252 13076 14254
rect 12908 14242 12964 14252
rect 12908 13860 12964 13870
rect 12572 13634 12628 13646
rect 12572 13582 12574 13634
rect 12626 13582 12628 13634
rect 12572 13522 12628 13582
rect 12908 13636 12964 13804
rect 12908 13542 12964 13580
rect 12572 13470 12574 13522
rect 12626 13470 12628 13522
rect 12572 13458 12628 13470
rect 12684 13076 12740 13086
rect 12684 13074 12964 13076
rect 12684 13022 12686 13074
rect 12738 13022 12964 13074
rect 12684 13020 12964 13022
rect 12684 13010 12740 13020
rect 12796 12850 12852 12862
rect 12796 12798 12798 12850
rect 12850 12798 12852 12850
rect 12796 12740 12852 12798
rect 12908 12850 12964 13020
rect 12908 12798 12910 12850
rect 12962 12798 12964 12850
rect 12908 12786 12964 12798
rect 12796 12674 12852 12684
rect 12908 12628 12964 12638
rect 12516 12460 12852 12516
rect 12236 12348 12404 12404
rect 12460 12384 12516 12460
rect 12796 12402 12852 12460
rect 11900 12290 11956 12302
rect 11900 12238 11902 12290
rect 11954 12238 11956 12290
rect 11788 11954 11844 11966
rect 11788 11902 11790 11954
rect 11842 11902 11844 11954
rect 11788 11732 11844 11902
rect 11788 11666 11844 11676
rect 11676 11554 11732 11564
rect 11788 11508 11844 11518
rect 11900 11508 11956 12238
rect 11788 11506 11956 11508
rect 11788 11454 11790 11506
rect 11842 11454 11956 11506
rect 11788 11452 11956 11454
rect 12012 12180 12068 12190
rect 12348 12180 12404 12348
rect 12796 12350 12798 12402
rect 12850 12350 12852 12402
rect 12796 12338 12852 12350
rect 11788 11442 11844 11452
rect 11676 11284 11732 11294
rect 11676 11190 11732 11228
rect 11900 11172 11956 11182
rect 11900 11078 11956 11116
rect 12012 10836 12068 12124
rect 12124 12124 12404 12180
rect 12572 12180 12628 12190
rect 12124 12066 12180 12124
rect 12124 12014 12126 12066
rect 12178 12014 12180 12066
rect 12124 12002 12180 12014
rect 12124 11396 12180 11406
rect 12124 11282 12180 11340
rect 12124 11230 12126 11282
rect 12178 11230 12180 11282
rect 12124 11218 12180 11230
rect 11788 10780 12068 10836
rect 11564 9996 11732 10052
rect 11116 9774 11118 9826
rect 11170 9774 11172 9826
rect 11116 9762 11172 9774
rect 11228 9772 11396 9828
rect 11564 9828 11620 9838
rect 10892 9716 10948 9726
rect 9660 8428 9828 8484
rect 9548 6402 9604 6412
rect 9660 8260 9716 8270
rect 9660 7364 9716 8204
rect 9660 6804 9716 7308
rect 9660 5124 9716 6748
rect 9772 6130 9828 8428
rect 9884 6804 9940 8652
rect 10332 8484 10388 8494
rect 9996 8370 10052 8382
rect 9996 8318 9998 8370
rect 10050 8318 10052 8370
rect 9996 7700 10052 8318
rect 9996 7634 10052 7644
rect 10332 7698 10388 8428
rect 10332 7646 10334 7698
rect 10386 7646 10388 7698
rect 10332 7634 10388 7646
rect 10556 7698 10612 8876
rect 10780 9268 10836 9278
rect 10668 8818 10724 8830
rect 10668 8766 10670 8818
rect 10722 8766 10724 8818
rect 10668 8260 10724 8766
rect 10668 8194 10724 8204
rect 10556 7646 10558 7698
rect 10610 7646 10612 7698
rect 10556 7634 10612 7646
rect 10108 7588 10164 7598
rect 10108 7494 10164 7532
rect 10668 7476 10724 7486
rect 10668 7382 10724 7420
rect 10220 7250 10276 7262
rect 10220 7198 10222 7250
rect 10274 7198 10276 7250
rect 9996 6804 10052 6814
rect 9884 6802 10052 6804
rect 9884 6750 9998 6802
rect 10050 6750 10052 6802
rect 9884 6748 10052 6750
rect 9884 6692 9940 6748
rect 9996 6738 10052 6748
rect 9884 6626 9940 6636
rect 9772 6078 9774 6130
rect 9826 6078 9828 6130
rect 9772 6066 9828 6078
rect 10220 5908 10276 7198
rect 10444 6468 10500 6478
rect 10332 6244 10388 6254
rect 10332 6130 10388 6188
rect 10332 6078 10334 6130
rect 10386 6078 10388 6130
rect 10332 6066 10388 6078
rect 10444 6130 10500 6412
rect 10444 6078 10446 6130
rect 10498 6078 10500 6130
rect 10444 6066 10500 6078
rect 9660 5122 9828 5124
rect 9660 5070 9662 5122
rect 9714 5070 9828 5122
rect 9660 5068 9828 5070
rect 9660 5058 9716 5068
rect 9212 4610 9268 4620
rect 9100 4498 9156 4508
rect 9772 4338 9828 5068
rect 10220 4788 10276 5852
rect 10332 5796 10388 5806
rect 10332 5234 10388 5740
rect 10556 5684 10612 5694
rect 10556 5590 10612 5628
rect 10332 5182 10334 5234
rect 10386 5182 10388 5234
rect 10332 5170 10388 5182
rect 10780 5010 10836 9212
rect 10892 9266 10948 9660
rect 10892 9214 10894 9266
rect 10946 9214 10948 9266
rect 10892 8372 10948 9214
rect 10892 8306 10948 8316
rect 11004 8818 11060 8830
rect 11004 8766 11006 8818
rect 11058 8766 11060 8818
rect 10780 4958 10782 5010
rect 10834 4958 10836 5010
rect 10780 4900 10836 4958
rect 10780 4834 10836 4844
rect 10892 4898 10948 4910
rect 10892 4846 10894 4898
rect 10946 4846 10948 4898
rect 10220 4722 10276 4732
rect 10892 4564 10948 4846
rect 10556 4508 10948 4564
rect 10556 4450 10612 4508
rect 10556 4398 10558 4450
rect 10610 4398 10612 4450
rect 10556 4386 10612 4398
rect 9772 4286 9774 4338
rect 9826 4286 9828 4338
rect 9772 4274 9828 4286
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 7868 3490 7924 3502
rect 8428 4226 8484 4238
rect 8428 4174 8430 4226
rect 8482 4174 8484 4226
rect 8428 3388 8484 4174
rect 10556 3666 10612 3678
rect 10556 3614 10558 3666
rect 10610 3614 10612 3666
rect 9772 3556 9828 3566
rect 9772 3462 9828 3500
rect 8092 3332 8484 3388
rect 8764 3442 8820 3454
rect 8764 3390 8766 3442
rect 8818 3390 8820 3442
rect 8764 3388 8820 3390
rect 8764 3332 9268 3388
rect 8092 980 8148 3332
rect 7868 924 8148 980
rect 7868 800 7924 924
rect 9212 800 9268 3332
rect 10556 800 10612 3614
rect 11004 3556 11060 8766
rect 11116 7252 11172 7262
rect 11116 6018 11172 7196
rect 11116 5966 11118 6018
rect 11170 5966 11172 6018
rect 11116 5954 11172 5966
rect 11116 5010 11172 5022
rect 11116 4958 11118 5010
rect 11170 4958 11172 5010
rect 11116 4452 11172 4958
rect 11228 4788 11284 9772
rect 11452 9602 11508 9614
rect 11452 9550 11454 9602
rect 11506 9550 11508 9602
rect 11452 8372 11508 9550
rect 11564 8820 11620 9772
rect 11564 8754 11620 8764
rect 11452 8306 11508 8316
rect 11676 8596 11732 9996
rect 11788 9826 11844 10780
rect 11788 9774 11790 9826
rect 11842 9774 11844 9826
rect 11788 9762 11844 9774
rect 11900 9940 11956 9950
rect 11900 9154 11956 9884
rect 11900 9102 11902 9154
rect 11954 9102 11956 9154
rect 11900 9090 11956 9102
rect 12012 9156 12068 9166
rect 11340 8260 11396 8270
rect 11340 6018 11396 8204
rect 11564 6132 11620 6142
rect 11564 6038 11620 6076
rect 11340 5966 11342 6018
rect 11394 5966 11396 6018
rect 11340 5954 11396 5966
rect 11676 6018 11732 8540
rect 11788 7364 11844 7374
rect 11788 7270 11844 7308
rect 12012 6020 12068 9100
rect 12124 8372 12180 8382
rect 12124 8278 12180 8316
rect 12236 8260 12292 12124
rect 12572 12086 12628 12124
rect 12908 12178 12964 12572
rect 12908 12126 12910 12178
rect 12962 12126 12964 12178
rect 12348 11844 12404 11854
rect 12348 10612 12404 11788
rect 12460 11732 12516 11742
rect 12460 10836 12516 11676
rect 12796 11732 12852 11742
rect 12796 11620 12852 11676
rect 12460 10770 12516 10780
rect 12572 11618 12852 11620
rect 12572 11566 12798 11618
rect 12850 11566 12852 11618
rect 12572 11564 12852 11566
rect 12348 10556 12516 10612
rect 12460 10052 12516 10556
rect 12236 8194 12292 8204
rect 12348 9996 12516 10052
rect 12572 10050 12628 11564
rect 12796 11554 12852 11564
rect 12908 11508 12964 12126
rect 12908 11442 12964 11452
rect 12572 9998 12574 10050
rect 12626 9998 12628 10050
rect 12236 7700 12292 7710
rect 12348 7700 12404 9996
rect 12572 9156 12628 9998
rect 12908 11284 12964 11294
rect 13020 11284 13076 14252
rect 13132 13860 13188 15092
rect 13580 14306 13636 14318
rect 13580 14254 13582 14306
rect 13634 14254 13636 14306
rect 13580 13972 13636 14254
rect 14140 14306 14196 14318
rect 14476 14308 14532 14318
rect 14140 14254 14142 14306
rect 14194 14254 14196 14306
rect 13580 13916 14084 13972
rect 13132 13794 13188 13804
rect 13356 13748 13412 13758
rect 13356 13654 13412 13692
rect 13692 13748 13748 13758
rect 13244 13522 13300 13534
rect 13244 13470 13246 13522
rect 13298 13470 13300 13522
rect 12908 11282 13076 11284
rect 12908 11230 12910 11282
rect 12962 11230 13076 11282
rect 12908 11228 13076 11230
rect 13132 12850 13188 12862
rect 13132 12798 13134 12850
rect 13186 12798 13188 12850
rect 12908 10724 12964 11228
rect 12796 9716 12852 9726
rect 12796 9622 12852 9660
rect 12572 9090 12628 9100
rect 12684 9602 12740 9614
rect 12684 9550 12686 9602
rect 12738 9550 12740 9602
rect 12292 7644 12404 7700
rect 12460 8260 12516 8270
rect 12124 6578 12180 6590
rect 12124 6526 12126 6578
rect 12178 6526 12180 6578
rect 12124 6132 12180 6526
rect 12124 6066 12180 6076
rect 11676 5966 11678 6018
rect 11730 5966 11732 6018
rect 11676 5954 11732 5966
rect 11900 5964 12068 6020
rect 11340 5012 11396 5022
rect 11340 4918 11396 4956
rect 11900 5010 11956 5964
rect 12236 5906 12292 7644
rect 12460 6018 12516 8204
rect 12460 5966 12462 6018
rect 12514 5966 12516 6018
rect 12460 5954 12516 5966
rect 12236 5854 12238 5906
rect 12290 5854 12292 5906
rect 12236 5842 12292 5854
rect 12124 5794 12180 5806
rect 12124 5742 12126 5794
rect 12178 5742 12180 5794
rect 11900 4958 11902 5010
rect 11954 4958 11956 5010
rect 11228 4722 11284 4732
rect 11116 4386 11172 4396
rect 11900 4452 11956 4958
rect 12012 5012 12068 5022
rect 12012 4918 12068 4956
rect 12124 4900 12180 5742
rect 12572 5124 12628 5134
rect 12572 5030 12628 5068
rect 12124 4806 12180 4844
rect 11900 4386 11956 4396
rect 12684 4452 12740 9550
rect 12796 8258 12852 8270
rect 12796 8206 12798 8258
rect 12850 8206 12852 8258
rect 12796 7364 12852 8206
rect 12796 6804 12852 7308
rect 12796 6690 12852 6748
rect 12796 6638 12798 6690
rect 12850 6638 12852 6690
rect 12796 6626 12852 6638
rect 12908 6468 12964 10668
rect 13020 10836 13076 10846
rect 13020 10722 13076 10780
rect 13020 10670 13022 10722
rect 13074 10670 13076 10722
rect 13020 10658 13076 10670
rect 13132 9828 13188 12798
rect 13244 12068 13300 13470
rect 13580 13522 13636 13534
rect 13580 13470 13582 13522
rect 13634 13470 13636 13522
rect 13468 12628 13524 12638
rect 13468 12290 13524 12572
rect 13468 12238 13470 12290
rect 13522 12238 13524 12290
rect 13468 12226 13524 12238
rect 13580 12290 13636 13470
rect 13692 12962 13748 13692
rect 13692 12910 13694 12962
rect 13746 12910 13748 12962
rect 13692 12898 13748 12910
rect 13916 13634 13972 13646
rect 13916 13582 13918 13634
rect 13970 13582 13972 13634
rect 13804 12740 13860 12750
rect 13804 12646 13860 12684
rect 13580 12238 13582 12290
rect 13634 12238 13636 12290
rect 13580 12180 13636 12238
rect 13580 12114 13636 12124
rect 13692 12628 13748 12638
rect 13244 12012 13412 12068
rect 13132 9762 13188 9772
rect 13244 11396 13300 11406
rect 12684 4386 12740 4396
rect 12796 6412 12964 6468
rect 13020 6692 13076 6702
rect 12684 4228 12740 4238
rect 12796 4228 12852 6412
rect 13020 6018 13076 6636
rect 13020 5966 13022 6018
rect 13074 5966 13076 6018
rect 13020 5954 13076 5966
rect 12684 4226 12852 4228
rect 12684 4174 12686 4226
rect 12738 4174 12852 4226
rect 12684 4172 12852 4174
rect 12908 5348 12964 5358
rect 12908 5234 12964 5292
rect 12908 5182 12910 5234
rect 12962 5182 12964 5234
rect 12908 4228 12964 5182
rect 13244 5124 13300 11340
rect 13356 11284 13412 12012
rect 13356 5908 13412 11228
rect 13580 11954 13636 11966
rect 13580 11902 13582 11954
rect 13634 11902 13636 11954
rect 13356 5842 13412 5852
rect 13468 7700 13524 7710
rect 13468 5684 13524 7644
rect 13580 6020 13636 11902
rect 13692 11956 13748 12572
rect 13916 12628 13972 13582
rect 14028 13300 14084 13916
rect 14140 13522 14196 14254
rect 14364 14306 14532 14308
rect 14364 14254 14478 14306
rect 14530 14254 14532 14306
rect 14364 14252 14532 14254
rect 14252 13860 14308 13870
rect 14252 13766 14308 13804
rect 14140 13470 14142 13522
rect 14194 13470 14196 13522
rect 14140 13458 14196 13470
rect 14028 13244 14196 13300
rect 13916 12562 13972 12572
rect 14028 12738 14084 12750
rect 14028 12686 14030 12738
rect 14082 12686 14084 12738
rect 13692 9938 13748 11900
rect 13692 9886 13694 9938
rect 13746 9886 13748 9938
rect 13692 9874 13748 9886
rect 13804 11732 13860 11742
rect 13804 10610 13860 11676
rect 13916 11508 13972 11518
rect 13916 11414 13972 11452
rect 13804 10558 13806 10610
rect 13858 10558 13860 10610
rect 13804 9940 13860 10558
rect 13804 9874 13860 9884
rect 13916 11172 13972 11182
rect 13916 9716 13972 11116
rect 13580 5954 13636 5964
rect 13804 9604 13860 9614
rect 13468 5618 13524 5628
rect 13244 5058 13300 5068
rect 13692 5572 13748 5582
rect 13580 4452 13636 4462
rect 12684 4162 12740 4172
rect 12908 4162 12964 4172
rect 13244 4226 13300 4238
rect 13244 4174 13246 4226
rect 13298 4174 13300 4226
rect 13244 4116 13300 4174
rect 13244 4050 13300 4060
rect 12236 3666 12292 3678
rect 12236 3614 12238 3666
rect 12290 3614 12292 3666
rect 11564 3556 11620 3566
rect 11004 3554 11620 3556
rect 11004 3502 11566 3554
rect 11618 3502 11620 3554
rect 11004 3500 11620 3502
rect 11564 3490 11620 3500
rect 12236 3388 12292 3614
rect 11900 3332 12292 3388
rect 13244 3668 13300 3678
rect 11900 800 11956 3332
rect 13244 800 13300 3612
rect 13580 3554 13636 4396
rect 13692 4338 13748 5516
rect 13804 5234 13860 9548
rect 13916 8146 13972 9660
rect 14028 8260 14084 12686
rect 14140 11284 14196 13244
rect 14364 12740 14420 14252
rect 14476 14242 14532 14252
rect 14700 13748 14756 13758
rect 14700 13634 14756 13692
rect 14700 13582 14702 13634
rect 14754 13582 14756 13634
rect 14588 13300 14644 13310
rect 14588 12964 14644 13244
rect 14364 12516 14420 12684
rect 14476 12850 14532 12862
rect 14476 12798 14478 12850
rect 14530 12798 14532 12850
rect 14476 12628 14532 12798
rect 14476 12562 14532 12572
rect 14588 12738 14644 12908
rect 14588 12686 14590 12738
rect 14642 12686 14644 12738
rect 14252 12460 14420 12516
rect 14252 12292 14308 12460
rect 14588 12404 14644 12686
rect 14252 12160 14308 12236
rect 14364 12348 14644 12404
rect 14364 12290 14420 12348
rect 14364 12238 14366 12290
rect 14418 12238 14420 12290
rect 14364 12226 14420 12238
rect 14476 12180 14532 12190
rect 14476 11396 14532 12124
rect 14140 11282 14308 11284
rect 14140 11230 14142 11282
rect 14194 11230 14308 11282
rect 14140 11228 14308 11230
rect 14140 11218 14196 11228
rect 14140 9716 14196 9726
rect 14140 8370 14196 9660
rect 14140 8318 14142 8370
rect 14194 8318 14196 8370
rect 14140 8306 14196 8318
rect 14028 8194 14084 8204
rect 13916 8094 13918 8146
rect 13970 8094 13972 8146
rect 13916 8082 13972 8094
rect 14028 8036 14084 8046
rect 14028 8034 14196 8036
rect 14028 7982 14030 8034
rect 14082 7982 14196 8034
rect 14028 7980 14196 7982
rect 14028 7970 14084 7980
rect 14028 7140 14084 7150
rect 13916 6804 13972 6814
rect 13916 6690 13972 6748
rect 13916 6638 13918 6690
rect 13970 6638 13972 6690
rect 13916 6626 13972 6638
rect 14028 6130 14084 7084
rect 14028 6078 14030 6130
rect 14082 6078 14084 6130
rect 14028 6066 14084 6078
rect 13804 5182 13806 5234
rect 13858 5182 13860 5234
rect 13804 5170 13860 5182
rect 13916 5684 13972 5694
rect 13692 4286 13694 4338
rect 13746 4286 13748 4338
rect 13692 4274 13748 4286
rect 13916 4338 13972 5628
rect 14028 5012 14084 5022
rect 14028 4564 14084 4956
rect 14028 4498 14084 4508
rect 13916 4286 13918 4338
rect 13970 4286 13972 4338
rect 13916 4274 13972 4286
rect 13580 3502 13582 3554
rect 13634 3502 13636 3554
rect 13580 3490 13636 3502
rect 14140 3556 14196 7980
rect 14252 7700 14308 11228
rect 14476 11172 14532 11340
rect 14476 11106 14532 11116
rect 14588 12178 14644 12190
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14252 7634 14308 7644
rect 14364 10610 14420 10622
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14252 6804 14308 6814
rect 14252 5122 14308 6748
rect 14252 5070 14254 5122
rect 14306 5070 14308 5122
rect 14252 5058 14308 5070
rect 14252 4564 14308 4574
rect 14364 4564 14420 10558
rect 14588 8258 14644 12126
rect 14700 11732 14756 13582
rect 14812 12628 14868 15092
rect 15036 14306 15092 15820
rect 15372 15874 15428 16270
rect 16268 16322 16324 16334
rect 16268 16270 16270 16322
rect 16322 16270 16324 16322
rect 16268 16210 16324 16270
rect 16268 16158 16270 16210
rect 16322 16158 16324 16210
rect 16268 16146 16324 16158
rect 15372 15822 15374 15874
rect 15426 15822 15428 15874
rect 15036 14254 15038 14306
rect 15090 14254 15092 14306
rect 14812 12562 14868 12572
rect 14924 13860 14980 13870
rect 14924 13636 14980 13804
rect 14700 11666 14756 11676
rect 14812 12404 14868 12414
rect 14812 11618 14868 12348
rect 14924 12292 14980 13580
rect 15036 12964 15092 14254
rect 15260 15202 15316 15214
rect 15260 15150 15262 15202
rect 15314 15150 15316 15202
rect 15260 14308 15316 15150
rect 15260 14242 15316 14252
rect 15148 14196 15204 14206
rect 15148 13970 15204 14140
rect 15148 13918 15150 13970
rect 15202 13918 15204 13970
rect 15148 13860 15204 13918
rect 15148 13794 15204 13804
rect 15092 12908 15316 12964
rect 15036 12898 15092 12908
rect 15148 12404 15204 12414
rect 15148 12310 15204 12348
rect 15036 12292 15092 12302
rect 14924 12290 15092 12292
rect 14924 12238 15038 12290
rect 15090 12238 15092 12290
rect 14924 12236 15092 12238
rect 15036 12180 15092 12236
rect 15036 12124 15204 12180
rect 14812 11566 14814 11618
rect 14866 11566 14868 11618
rect 14812 11554 14868 11566
rect 14700 11284 14756 11294
rect 14700 11190 14756 11228
rect 14700 10724 14756 10734
rect 14700 10722 14980 10724
rect 14700 10670 14702 10722
rect 14754 10670 14980 10722
rect 14700 10668 14980 10670
rect 14700 10658 14756 10668
rect 14588 8206 14590 8258
rect 14642 8206 14644 8258
rect 14588 8194 14644 8206
rect 14812 8260 14868 8270
rect 14700 6578 14756 6590
rect 14700 6526 14702 6578
rect 14754 6526 14756 6578
rect 14700 6130 14756 6526
rect 14700 6078 14702 6130
rect 14754 6078 14756 6130
rect 14700 6066 14756 6078
rect 14812 6018 14868 8204
rect 14812 5966 14814 6018
rect 14866 5966 14868 6018
rect 14812 5954 14868 5966
rect 14476 5908 14532 5918
rect 14476 5814 14532 5852
rect 14252 4562 14420 4564
rect 14252 4510 14254 4562
rect 14306 4510 14420 4562
rect 14252 4508 14420 4510
rect 14252 4498 14308 4508
rect 14924 4338 14980 10668
rect 15148 8708 15204 12124
rect 15260 11844 15316 12908
rect 15372 12404 15428 15822
rect 15708 15876 15764 15886
rect 15708 15540 15764 15820
rect 15708 15474 15764 15484
rect 16044 15876 16100 15886
rect 15820 15204 15876 15214
rect 15820 15092 15988 15148
rect 15820 15072 15876 15092
rect 15484 14420 15540 14430
rect 15484 13972 15540 14364
rect 15596 14308 15652 14318
rect 15652 14252 15764 14308
rect 15596 14176 15652 14252
rect 15596 13972 15652 13982
rect 15484 13970 15652 13972
rect 15484 13918 15598 13970
rect 15650 13918 15652 13970
rect 15484 13916 15652 13918
rect 15596 13906 15652 13916
rect 15708 13636 15764 14252
rect 15708 13570 15764 13580
rect 15932 12964 15988 15092
rect 16044 14308 16100 15820
rect 16716 15874 16772 15886
rect 16716 15822 16718 15874
rect 16770 15822 16772 15874
rect 16716 15428 16772 15822
rect 17164 15874 17220 15886
rect 17164 15822 17166 15874
rect 17218 15822 17220 15874
rect 16716 15372 17108 15428
rect 16492 15204 16548 15214
rect 16940 15204 16996 15214
rect 16492 15202 16996 15204
rect 16492 15150 16494 15202
rect 16546 15150 16942 15202
rect 16994 15150 16996 15202
rect 16492 15148 16996 15150
rect 16492 15138 16548 15148
rect 16604 14868 16660 14878
rect 16492 14644 16548 14654
rect 16044 14306 16212 14308
rect 16044 14254 16046 14306
rect 16098 14254 16212 14306
rect 16044 14252 16212 14254
rect 16044 14242 16100 14252
rect 16044 13636 16100 13646
rect 16044 13542 16100 13580
rect 16156 13522 16212 14252
rect 16156 13470 16158 13522
rect 16210 13470 16212 13522
rect 16156 13458 16212 13470
rect 16492 14306 16548 14588
rect 16492 14254 16494 14306
rect 16546 14254 16548 14306
rect 15932 12908 16212 12964
rect 15484 12738 15540 12750
rect 15484 12686 15486 12738
rect 15538 12686 15540 12738
rect 15484 12628 15540 12686
rect 15484 12562 15540 12572
rect 15932 12738 15988 12750
rect 15932 12686 15934 12738
rect 15986 12686 15988 12738
rect 15820 12404 15876 12414
rect 15372 12348 15652 12404
rect 15372 12180 15428 12190
rect 15372 12178 15540 12180
rect 15372 12126 15374 12178
rect 15426 12126 15540 12178
rect 15372 12124 15540 12126
rect 15372 12114 15428 12124
rect 15260 11778 15316 11788
rect 15372 11170 15428 11182
rect 15372 11118 15374 11170
rect 15426 11118 15428 11170
rect 15372 11060 15428 11118
rect 15372 10994 15428 11004
rect 15484 10498 15540 12124
rect 15596 11956 15652 12348
rect 15820 12068 15876 12348
rect 15820 12002 15876 12012
rect 15596 11890 15652 11900
rect 15820 11844 15876 11854
rect 15484 10446 15486 10498
rect 15538 10446 15540 10498
rect 15148 8652 15428 8708
rect 15260 8484 15316 8494
rect 15148 8372 15204 8382
rect 15148 8278 15204 8316
rect 15036 8260 15092 8270
rect 15036 8166 15092 8204
rect 15260 8258 15316 8428
rect 15260 8206 15262 8258
rect 15314 8206 15316 8258
rect 15260 8194 15316 8206
rect 15372 6692 15428 8652
rect 15036 5908 15092 5918
rect 15036 5814 15092 5852
rect 15372 5684 15428 6636
rect 15484 5906 15540 10446
rect 15596 11732 15652 11742
rect 15596 8484 15652 11676
rect 15820 10500 15876 11788
rect 15932 11620 15988 12686
rect 15932 11554 15988 11564
rect 16044 11844 16100 11854
rect 15932 11396 15988 11406
rect 15932 11302 15988 11340
rect 15820 10498 15988 10500
rect 15820 10446 15822 10498
rect 15874 10446 15988 10498
rect 15820 10444 15988 10446
rect 15820 10434 15876 10444
rect 15820 9716 15876 9726
rect 15596 8418 15652 8428
rect 15708 9714 15876 9716
rect 15708 9662 15822 9714
rect 15874 9662 15876 9714
rect 15708 9660 15876 9662
rect 15708 8372 15764 9660
rect 15820 9650 15876 9660
rect 15932 9492 15988 10444
rect 15708 8306 15764 8316
rect 15820 9436 15988 9492
rect 15484 5854 15486 5906
rect 15538 5854 15540 5906
rect 15484 5842 15540 5854
rect 15820 5908 15876 9436
rect 16044 7924 16100 11788
rect 15932 6020 15988 6030
rect 16044 6020 16100 7868
rect 16156 9828 16212 12908
rect 16268 12740 16324 12750
rect 16268 12646 16324 12684
rect 16380 12404 16436 12414
rect 16492 12404 16548 14254
rect 16604 13970 16660 14812
rect 16604 13918 16606 13970
rect 16658 13918 16660 13970
rect 16604 13906 16660 13918
rect 16380 12402 16548 12404
rect 16380 12350 16382 12402
rect 16434 12350 16548 12402
rect 16380 12348 16548 12350
rect 16604 13522 16660 13534
rect 16604 13470 16606 13522
rect 16658 13470 16660 13522
rect 16380 12338 16436 12348
rect 16604 12292 16660 13470
rect 16492 12236 16660 12292
rect 16492 10724 16548 12236
rect 16716 11732 16772 15148
rect 16940 15138 16996 15148
rect 16940 14754 16996 14766
rect 16940 14702 16942 14754
rect 16994 14702 16996 14754
rect 16940 14308 16996 14702
rect 16828 14306 16996 14308
rect 16828 14254 16942 14306
rect 16994 14254 16996 14306
rect 16828 14252 16996 14254
rect 16828 13748 16884 14252
rect 16940 14242 16996 14252
rect 17052 14308 17108 15372
rect 17052 14242 17108 14252
rect 17164 14196 17220 15822
rect 17276 14754 17332 17164
rect 17612 16884 17668 16894
rect 17612 16790 17668 16828
rect 17612 15876 17668 15886
rect 17500 15874 17668 15876
rect 17500 15822 17614 15874
rect 17666 15822 17668 15874
rect 17500 15820 17668 15822
rect 17500 15092 17556 15820
rect 17612 15810 17668 15820
rect 17948 15876 18004 15886
rect 17948 15782 18004 15820
rect 18172 15540 18228 18508
rect 18284 16884 18340 16894
rect 18284 16790 18340 16828
rect 18284 15540 18340 15550
rect 18172 15538 18340 15540
rect 18172 15486 18286 15538
rect 18338 15486 18340 15538
rect 18172 15484 18340 15486
rect 17836 15204 17892 15214
rect 17500 15026 17556 15036
rect 17612 15202 17892 15204
rect 17612 15150 17838 15202
rect 17890 15150 17892 15202
rect 17612 15148 17892 15150
rect 17276 14702 17278 14754
rect 17330 14702 17332 14754
rect 17276 14690 17332 14702
rect 17164 14130 17220 14140
rect 17388 14308 17444 14318
rect 16940 13972 16996 13982
rect 16940 13878 16996 13916
rect 17388 13748 17444 14252
rect 16828 13692 16996 13748
rect 16828 12738 16884 12750
rect 16828 12686 16830 12738
rect 16882 12686 16884 12738
rect 16828 12292 16884 12686
rect 16828 12226 16884 12236
rect 16940 12180 16996 13692
rect 17388 13682 17444 13692
rect 17612 13636 17668 15148
rect 17836 15138 17892 15148
rect 18172 14644 18228 15484
rect 18284 15474 18340 15484
rect 18060 14588 18172 14644
rect 17948 14532 18004 14542
rect 17948 13972 18004 14476
rect 17276 12852 17332 12862
rect 17276 12758 17332 12796
rect 16940 12114 16996 12124
rect 16492 10386 16548 10668
rect 16604 11508 16660 11518
rect 16604 11394 16660 11452
rect 16604 11342 16606 11394
rect 16658 11342 16660 11394
rect 16604 10612 16660 11342
rect 16604 10546 16660 10556
rect 16492 10334 16494 10386
rect 16546 10334 16548 10386
rect 16492 10164 16548 10334
rect 16604 10388 16660 10398
rect 16604 10294 16660 10332
rect 16492 10108 16660 10164
rect 16492 9828 16548 9838
rect 16156 9826 16548 9828
rect 16156 9774 16494 9826
rect 16546 9774 16548 9826
rect 16156 9772 16548 9774
rect 16156 8258 16212 9772
rect 16492 9762 16548 9772
rect 16156 8206 16158 8258
rect 16210 8206 16212 8258
rect 16156 6804 16212 8206
rect 16604 7252 16660 10108
rect 16716 9042 16772 11676
rect 16828 12066 16884 12078
rect 16828 12014 16830 12066
rect 16882 12014 16884 12066
rect 16828 11508 16884 12014
rect 17612 12066 17668 13580
rect 17836 13748 17892 13758
rect 17836 12850 17892 13692
rect 17948 13746 18004 13916
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13682 18004 13694
rect 17836 12798 17838 12850
rect 17890 12798 17892 12850
rect 17612 12014 17614 12066
rect 17666 12014 17668 12066
rect 16940 11956 16996 11966
rect 16940 11954 17556 11956
rect 16940 11902 16942 11954
rect 16994 11902 17556 11954
rect 16940 11900 17556 11902
rect 16940 11890 16996 11900
rect 16828 11452 17108 11508
rect 16940 11284 16996 11294
rect 16828 11172 16884 11182
rect 16828 10610 16884 11116
rect 16940 10722 16996 11228
rect 16940 10670 16942 10722
rect 16994 10670 16996 10722
rect 16940 10658 16996 10670
rect 16828 10558 16830 10610
rect 16882 10558 16884 10610
rect 16828 10546 16884 10558
rect 17052 9156 17108 11452
rect 17276 11284 17332 11294
rect 17276 11190 17332 11228
rect 17500 10500 17556 11900
rect 17612 11954 17668 12014
rect 17612 11902 17614 11954
rect 17666 11902 17668 11954
rect 17612 11890 17668 11902
rect 17724 12738 17780 12750
rect 17724 12686 17726 12738
rect 17778 12686 17780 12738
rect 17724 11844 17780 12686
rect 17724 11778 17780 11788
rect 17836 11060 17892 12798
rect 17724 11004 17892 11060
rect 17948 11954 18004 11966
rect 17948 11902 17950 11954
rect 18002 11902 18004 11954
rect 17500 10434 17556 10444
rect 17612 10724 17668 10734
rect 17612 10050 17668 10668
rect 17724 10276 17780 11004
rect 17948 10948 18004 11902
rect 17948 10834 18004 10892
rect 17948 10782 17950 10834
rect 18002 10782 18004 10834
rect 17948 10770 18004 10782
rect 17724 10210 17780 10220
rect 17948 10498 18004 10510
rect 17948 10446 17950 10498
rect 18002 10446 18004 10498
rect 17612 9998 17614 10050
rect 17666 9998 17668 10050
rect 17612 9986 17668 9998
rect 17724 10052 17780 10062
rect 17276 9826 17332 9838
rect 17276 9774 17278 9826
rect 17330 9774 17332 9826
rect 17052 9090 17108 9100
rect 17164 9714 17220 9726
rect 17164 9662 17166 9714
rect 17218 9662 17220 9714
rect 16716 8990 16718 9042
rect 16770 8990 16772 9042
rect 16716 7474 16772 8990
rect 16828 8372 16884 8382
rect 17164 8372 17220 9662
rect 17276 8932 17332 9774
rect 17500 9828 17556 9866
rect 17500 9762 17556 9772
rect 17724 9716 17780 9996
rect 17724 9650 17780 9660
rect 17276 8866 17332 8876
rect 17612 9380 17668 9390
rect 16828 8370 17220 8372
rect 16828 8318 16830 8370
rect 16882 8318 17220 8370
rect 16828 8316 17220 8318
rect 17388 8708 17444 8718
rect 16828 8306 16884 8316
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16716 7410 16772 7422
rect 16604 7196 16772 7252
rect 16156 6738 16212 6748
rect 16604 7028 16660 7038
rect 16604 6130 16660 6972
rect 16604 6078 16606 6130
rect 16658 6078 16660 6130
rect 16604 6066 16660 6078
rect 16716 6580 16772 7196
rect 17276 6916 17332 6926
rect 17276 6822 17332 6860
rect 16716 6132 16772 6524
rect 16828 6802 16884 6814
rect 16828 6750 16830 6802
rect 16882 6750 16884 6802
rect 16828 6692 16884 6750
rect 16828 6356 16884 6636
rect 16828 6290 16884 6300
rect 17052 6692 17108 6702
rect 16828 6132 16884 6142
rect 16716 6076 16828 6132
rect 15932 6018 16100 6020
rect 15932 5966 15934 6018
rect 15986 5966 16100 6018
rect 15932 5964 16100 5966
rect 16156 6020 16212 6030
rect 15932 5954 15988 5964
rect 16156 5926 16212 5964
rect 15820 5842 15876 5852
rect 15372 5618 15428 5628
rect 15708 5794 15764 5806
rect 15708 5742 15710 5794
rect 15762 5742 15764 5794
rect 15036 5236 15092 5246
rect 15036 5142 15092 5180
rect 15708 5236 15764 5742
rect 15708 5170 15764 5180
rect 14924 4286 14926 4338
rect 14978 4286 14980 4338
rect 14924 4274 14980 4286
rect 15596 4676 15652 4686
rect 14588 4228 14644 4238
rect 14252 3668 14308 3678
rect 14252 3574 14308 3612
rect 14140 3490 14196 3500
rect 14588 800 14644 4172
rect 15484 4228 15540 4238
rect 15484 4134 15540 4172
rect 15596 3554 15652 4620
rect 16604 4452 16660 4462
rect 16716 4452 16772 6076
rect 16828 6038 16884 6076
rect 16940 6020 16996 6030
rect 16940 5926 16996 5964
rect 16828 5460 16884 5470
rect 16828 4562 16884 5404
rect 16828 4510 16830 4562
rect 16882 4510 16884 4562
rect 16828 4498 16884 4510
rect 16604 4450 16772 4452
rect 16604 4398 16606 4450
rect 16658 4398 16772 4450
rect 16604 4396 16772 4398
rect 16604 4386 16660 4396
rect 16940 4228 16996 4238
rect 17052 4228 17108 6636
rect 17388 6578 17444 8652
rect 17388 6526 17390 6578
rect 17442 6526 17444 6578
rect 17388 6514 17444 6526
rect 17612 6466 17668 9324
rect 17724 9268 17780 9278
rect 17724 9174 17780 9212
rect 17948 8708 18004 10446
rect 17948 8642 18004 8652
rect 18060 8372 18116 14588
rect 18172 14578 18228 14588
rect 18172 14306 18228 14318
rect 18172 14254 18174 14306
rect 18226 14254 18228 14306
rect 18172 12180 18228 14254
rect 18396 13524 18452 39004
rect 21980 39060 22036 43200
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 21980 38994 22036 39004
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 30044 27076 30100 27086
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 27020 24612 27076 24622
rect 25228 23940 25284 23950
rect 24780 23828 24836 23838
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 23324 22484 23380 22494
rect 18620 22148 18676 22158
rect 18620 17778 18676 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 21644 21924 21700 21934
rect 19628 21252 19684 21262
rect 18620 17726 18622 17778
rect 18674 17726 18676 17778
rect 18620 17714 18676 17726
rect 19068 18004 19124 18014
rect 19068 17778 19124 17948
rect 19068 17726 19070 17778
rect 19122 17726 19124 17778
rect 19068 17714 19124 17726
rect 19516 17444 19572 17454
rect 19404 17442 19572 17444
rect 19404 17390 19518 17442
rect 19570 17390 19572 17442
rect 19404 17388 19572 17390
rect 18732 17108 18788 17118
rect 18732 17014 18788 17052
rect 18396 13458 18452 13468
rect 18508 16884 18564 16894
rect 18508 13076 18564 16828
rect 19068 16772 19124 16782
rect 19068 16678 19124 16716
rect 18732 16324 18788 16334
rect 18732 16210 18788 16268
rect 19180 16212 19236 16222
rect 18732 16158 18734 16210
rect 18786 16158 18788 16210
rect 18620 14980 18676 14990
rect 18620 14642 18676 14924
rect 18620 14590 18622 14642
rect 18674 14590 18676 14642
rect 18620 14578 18676 14590
rect 18620 13636 18676 13646
rect 18620 13542 18676 13580
rect 18508 13020 18676 13076
rect 18508 12850 18564 12862
rect 18508 12798 18510 12850
rect 18562 12798 18564 12850
rect 18172 12114 18228 12124
rect 18396 12738 18452 12750
rect 18396 12686 18398 12738
rect 18450 12686 18452 12738
rect 18284 12068 18340 12078
rect 18284 11974 18340 12012
rect 18172 11954 18228 11966
rect 18172 11902 18174 11954
rect 18226 11902 18228 11954
rect 18172 10724 18228 11902
rect 18172 10592 18228 10668
rect 18284 10836 18340 10846
rect 18172 10388 18228 10398
rect 18172 9268 18228 10332
rect 18284 9826 18340 10780
rect 18396 10052 18452 12686
rect 18396 9986 18452 9996
rect 18284 9774 18286 9826
rect 18338 9774 18340 9826
rect 18284 9492 18340 9774
rect 18284 9426 18340 9436
rect 18396 9604 18452 9614
rect 18284 9268 18340 9278
rect 18172 9266 18340 9268
rect 18172 9214 18286 9266
rect 18338 9214 18340 9266
rect 18172 9212 18340 9214
rect 18284 9202 18340 9212
rect 18172 8932 18228 8942
rect 18172 8838 18228 8876
rect 18396 8484 18452 9548
rect 18508 9380 18564 12798
rect 18620 9828 18676 13020
rect 18732 12628 18788 16158
rect 18956 16156 19180 16212
rect 18844 15202 18900 15214
rect 18844 15150 18846 15202
rect 18898 15150 18900 15202
rect 18844 14308 18900 15150
rect 18844 14242 18900 14252
rect 18732 10836 18788 12572
rect 18844 12740 18900 12750
rect 18844 12292 18900 12684
rect 18956 12516 19012 16156
rect 19180 16118 19236 16156
rect 19180 15202 19236 15214
rect 19180 15150 19182 15202
rect 19234 15150 19236 15202
rect 19068 14306 19124 14318
rect 19068 14254 19070 14306
rect 19122 14254 19124 14306
rect 19068 14084 19124 14254
rect 19068 14018 19124 14028
rect 19180 13748 19236 15150
rect 19180 13682 19236 13692
rect 19404 13188 19460 17388
rect 19516 17378 19572 17388
rect 19516 17220 19572 17230
rect 19516 17106 19572 17164
rect 19516 17054 19518 17106
rect 19570 17054 19572 17106
rect 19516 16996 19572 17054
rect 19516 16930 19572 16940
rect 19628 16212 19684 21196
rect 21084 20580 21140 20590
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20244 20356 20254
rect 20300 20132 20580 20188
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18564 19908 18574
rect 19852 17778 19908 18508
rect 20076 18340 20132 18350
rect 20076 18246 20132 18284
rect 19852 17726 19854 17778
rect 19906 17726 19908 17778
rect 19852 17714 19908 17726
rect 20412 17444 20468 17454
rect 20300 17442 20468 17444
rect 20300 17390 20414 17442
rect 20466 17390 20468 17442
rect 20300 17388 20468 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17220 20244 17230
rect 19964 17108 20020 17118
rect 20188 17108 20244 17164
rect 19964 17106 20244 17108
rect 19964 17054 19966 17106
rect 20018 17054 20244 17106
rect 19964 17052 20244 17054
rect 19964 17042 20020 17052
rect 19516 16156 19684 16212
rect 20188 16660 20244 16670
rect 19516 14420 19572 16156
rect 19740 15876 19796 15886
rect 19628 15874 19796 15876
rect 19628 15822 19742 15874
rect 19794 15822 19796 15874
rect 19628 15820 19796 15822
rect 19628 14532 19684 15820
rect 19740 15810 19796 15820
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19964 15540 20020 15550
rect 20188 15540 20244 16604
rect 20020 15484 20244 15540
rect 19964 15446 20020 15484
rect 19628 14466 19684 14476
rect 20076 14980 20132 14990
rect 20076 14530 20132 14924
rect 20076 14478 20078 14530
rect 20130 14478 20132 14530
rect 20076 14466 20132 14478
rect 19516 14354 19572 14364
rect 20188 14418 20244 15484
rect 20188 14366 20190 14418
rect 20242 14366 20244 14418
rect 20188 14354 20244 14366
rect 19628 14306 19684 14318
rect 19628 14254 19630 14306
rect 19682 14254 19684 14306
rect 19628 13972 19684 14254
rect 20188 14196 20244 14206
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13906 19684 13916
rect 19404 13122 19460 13132
rect 19740 13748 19796 13758
rect 19068 12964 19124 12974
rect 19068 12962 19572 12964
rect 19068 12910 19070 12962
rect 19122 12910 19572 12962
rect 19068 12908 19572 12910
rect 19068 12898 19124 12908
rect 19404 12740 19460 12750
rect 19292 12738 19460 12740
rect 19292 12686 19406 12738
rect 19458 12686 19460 12738
rect 19292 12684 19460 12686
rect 18956 12460 19124 12516
rect 18844 12198 18900 12236
rect 18956 12290 19012 12302
rect 18956 12238 18958 12290
rect 19010 12238 19012 12290
rect 18956 12180 19012 12238
rect 18956 12114 19012 12124
rect 18732 10770 18788 10780
rect 18844 11396 18900 11406
rect 18844 10722 18900 11340
rect 19068 10948 19124 12460
rect 18844 10670 18846 10722
rect 18898 10670 18900 10722
rect 18732 10388 18788 10398
rect 18732 10294 18788 10332
rect 18620 9772 18788 9828
rect 18620 9604 18676 9614
rect 18620 9510 18676 9548
rect 18508 9324 18676 9380
rect 18508 9156 18564 9166
rect 18508 9062 18564 9100
rect 18396 8418 18452 8428
rect 17836 7476 17892 7486
rect 18060 7476 18116 8316
rect 17836 7474 18116 7476
rect 17836 7422 17838 7474
rect 17890 7422 18116 7474
rect 17836 7420 18116 7422
rect 17836 7410 17892 7420
rect 18508 7362 18564 7374
rect 18508 7310 18510 7362
rect 18562 7310 18564 7362
rect 18284 7028 18340 7038
rect 17612 6414 17614 6466
rect 17666 6414 17668 6466
rect 17612 6356 17668 6414
rect 17164 6300 17668 6356
rect 17164 5234 17220 6300
rect 17612 6020 17668 6300
rect 17612 5954 17668 5964
rect 17724 6580 17780 6590
rect 17164 5182 17166 5234
rect 17218 5182 17220 5234
rect 17164 4340 17220 5182
rect 17164 4274 17220 4284
rect 17276 5236 17332 5246
rect 16940 4226 17108 4228
rect 16940 4174 16942 4226
rect 16994 4174 17108 4226
rect 16940 4172 17108 4174
rect 16940 4162 16996 4172
rect 15596 3502 15598 3554
rect 15650 3502 15652 3554
rect 15596 3490 15652 3502
rect 16156 3666 16212 3678
rect 16156 3614 16158 3666
rect 16210 3614 16212 3666
rect 16156 3388 16212 3614
rect 15932 3332 16212 3388
rect 15932 800 15988 3332
rect 17276 800 17332 5180
rect 17724 5122 17780 6524
rect 17836 6578 17892 6590
rect 17836 6526 17838 6578
rect 17890 6526 17892 6578
rect 17836 6356 17892 6526
rect 17836 6290 17892 6300
rect 18284 6132 18340 6972
rect 18508 6692 18564 7310
rect 18508 6626 18564 6636
rect 18620 7364 18676 9324
rect 18620 6690 18676 7308
rect 18620 6638 18622 6690
rect 18674 6638 18676 6690
rect 18396 6468 18452 6478
rect 18396 6374 18452 6412
rect 18508 6466 18564 6478
rect 18508 6414 18510 6466
rect 18562 6414 18564 6466
rect 18284 6066 18340 6076
rect 17724 5070 17726 5122
rect 17778 5070 17780 5122
rect 17724 5058 17780 5070
rect 17836 6018 17892 6030
rect 17836 5966 17838 6018
rect 17890 5966 17892 6018
rect 17836 4226 17892 5966
rect 17948 5908 18004 5918
rect 17948 5814 18004 5852
rect 18508 5460 18564 6414
rect 18620 5906 18676 6638
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5842 18676 5854
rect 18508 5394 18564 5404
rect 18396 5236 18452 5246
rect 18396 5142 18452 5180
rect 18732 5012 18788 9772
rect 18844 9716 18900 10670
rect 18844 9650 18900 9660
rect 18956 10892 19124 10948
rect 19180 12178 19236 12190
rect 19180 12126 19182 12178
rect 19234 12126 19236 12178
rect 18956 9380 19012 10892
rect 19068 10724 19124 10734
rect 19068 10630 19124 10668
rect 19180 10052 19236 12126
rect 19180 9986 19236 9996
rect 19068 9828 19124 9838
rect 19068 9734 19124 9772
rect 19180 9826 19236 9838
rect 19180 9774 19182 9826
rect 19234 9774 19236 9826
rect 18844 9324 19012 9380
rect 19180 9716 19236 9774
rect 18844 8932 18900 9324
rect 18844 8866 18900 8876
rect 18956 9156 19012 9166
rect 19180 9156 19236 9660
rect 18956 8370 19012 9100
rect 18956 8318 18958 8370
rect 19010 8318 19012 8370
rect 18956 8306 19012 8318
rect 19068 9100 19236 9156
rect 18956 6692 19012 6702
rect 19068 6692 19124 9100
rect 19180 8932 19236 8970
rect 19180 8866 19236 8876
rect 18956 6690 19124 6692
rect 18956 6638 18958 6690
rect 19010 6638 19124 6690
rect 18956 6636 19124 6638
rect 19180 8708 19236 8718
rect 18956 5682 19012 6636
rect 19068 6020 19124 6030
rect 19068 5906 19124 5964
rect 19068 5854 19070 5906
rect 19122 5854 19124 5906
rect 19068 5842 19124 5854
rect 18956 5630 18958 5682
rect 19010 5630 19012 5682
rect 18956 5618 19012 5630
rect 18732 4452 18788 4956
rect 18732 4386 18788 4396
rect 17836 4174 17838 4226
rect 17890 4174 17892 4226
rect 17836 3668 17892 4174
rect 17836 3602 17892 3612
rect 18620 3666 18676 3678
rect 18620 3614 18622 3666
rect 18674 3614 18676 3666
rect 17612 3556 17668 3566
rect 17612 3462 17668 3500
rect 18620 800 18676 3614
rect 19180 3556 19236 8652
rect 19292 6692 19348 12684
rect 19404 12674 19460 12684
rect 19404 12068 19460 12078
rect 19404 11506 19460 12012
rect 19404 11454 19406 11506
rect 19458 11454 19460 11506
rect 19404 11442 19460 11454
rect 19516 11508 19572 12908
rect 19740 12962 19796 13692
rect 19740 12910 19742 12962
rect 19794 12910 19796 12962
rect 19740 12898 19796 12910
rect 19628 12738 19684 12750
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19628 11956 19684 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 11890 19684 11900
rect 20188 11844 20244 14140
rect 20188 11778 20244 11788
rect 19516 10948 19572 11452
rect 19964 11396 20020 11406
rect 19964 11302 20020 11340
rect 20188 11394 20244 11406
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19516 10882 19572 10892
rect 20076 10836 20132 10846
rect 19516 10724 19572 10734
rect 19516 10050 19572 10668
rect 19964 10612 20020 10622
rect 19964 10518 20020 10556
rect 19516 9998 19518 10050
rect 19570 9998 19572 10050
rect 19516 9986 19572 9998
rect 19404 9940 19460 9950
rect 19404 8708 19460 9884
rect 20076 9604 20132 10780
rect 20188 10724 20244 11342
rect 20188 10658 20244 10668
rect 20076 9548 20244 9604
rect 19516 9492 19572 9502
rect 19516 9044 19572 9436
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9548
rect 19516 8932 19572 8988
rect 19964 9212 20244 9268
rect 19628 8932 19684 8942
rect 19516 8930 19684 8932
rect 19516 8878 19630 8930
rect 19682 8878 19684 8930
rect 19516 8876 19684 8878
rect 19628 8866 19684 8876
rect 19404 8652 19684 8708
rect 19628 8482 19684 8652
rect 19628 8430 19630 8482
rect 19682 8430 19684 8482
rect 19628 8418 19684 8430
rect 19964 8260 20020 9212
rect 19964 8128 20020 8204
rect 19740 8036 19796 8074
rect 19740 7970 19796 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19852 7700 19908 7710
rect 20300 7700 20356 17388
rect 20412 17378 20468 17388
rect 20412 16884 20468 16894
rect 20524 16884 20580 20132
rect 20972 19796 21028 19806
rect 20748 19684 20804 19694
rect 20412 16882 20580 16884
rect 20412 16830 20414 16882
rect 20466 16830 20580 16882
rect 20412 16828 20580 16830
rect 20412 16818 20468 16828
rect 20412 16324 20468 16334
rect 20412 16210 20468 16268
rect 20412 16158 20414 16210
rect 20466 16158 20468 16210
rect 20412 16146 20468 16158
rect 20524 14420 20580 16828
rect 20636 18450 20692 18462
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20636 15314 20692 18398
rect 20748 16322 20804 19628
rect 20860 19010 20916 19022
rect 20860 18958 20862 19010
rect 20914 18958 20916 19010
rect 20860 18452 20916 18958
rect 20860 18386 20916 18396
rect 20860 17780 20916 17790
rect 20860 17686 20916 17724
rect 20748 16270 20750 16322
rect 20802 16270 20804 16322
rect 20748 16258 20804 16270
rect 20860 16884 20916 16894
rect 20972 16884 21028 19740
rect 20860 16882 21028 16884
rect 20860 16830 20862 16882
rect 20914 16830 21028 16882
rect 20860 16828 21028 16830
rect 21084 17220 21140 20524
rect 21644 19346 21700 21868
rect 22988 21364 23044 21374
rect 22988 20914 23044 21308
rect 22988 20862 22990 20914
rect 23042 20862 23044 20914
rect 22988 20850 23044 20862
rect 22876 20804 22932 20814
rect 22876 20244 22932 20748
rect 23324 20188 23380 22428
rect 24780 22482 24836 23772
rect 24780 22430 24782 22482
rect 24834 22430 24836 22482
rect 24780 22148 24836 22430
rect 25228 22482 25284 23884
rect 26012 23604 26068 23614
rect 25228 22430 25230 22482
rect 25282 22430 25284 22482
rect 25228 22418 25284 22430
rect 25564 23044 25620 23054
rect 25564 22484 25620 22988
rect 26012 22484 26068 23548
rect 26460 23156 26516 23166
rect 25564 22352 25620 22428
rect 25900 22482 26068 22484
rect 25900 22430 26014 22482
rect 26066 22430 26068 22482
rect 25900 22428 26068 22430
rect 24780 22082 24836 22092
rect 25564 22260 25620 22270
rect 24108 21474 24164 21486
rect 24108 21422 24110 21474
rect 24162 21422 24164 21474
rect 24108 21364 24164 21422
rect 24556 21476 24612 21486
rect 24556 21382 24612 21420
rect 24892 21474 24948 21486
rect 24892 21422 24894 21474
rect 24946 21422 24948 21474
rect 24108 21298 24164 21308
rect 23436 21140 23492 21150
rect 23436 20914 23492 21084
rect 23436 20862 23438 20914
rect 23490 20862 23492 20914
rect 23436 20850 23492 20862
rect 23884 20916 23940 20926
rect 23884 20822 23940 20860
rect 24332 20692 24388 20702
rect 24332 20598 24388 20636
rect 24668 20580 24724 20590
rect 24668 20486 24724 20524
rect 22876 20130 22932 20188
rect 22876 20078 22878 20130
rect 22930 20078 22932 20130
rect 22876 20066 22932 20078
rect 23212 20132 23380 20188
rect 24892 20188 24948 21422
rect 25564 21476 25620 22204
rect 25564 21382 25620 21420
rect 25228 20578 25284 20590
rect 25228 20526 25230 20578
rect 25282 20526 25284 20578
rect 25228 20188 25284 20526
rect 25788 20578 25844 20590
rect 25788 20526 25790 20578
rect 25842 20526 25844 20578
rect 25788 20468 25844 20526
rect 25788 20188 25844 20412
rect 24892 20132 25172 20188
rect 25228 20132 25396 20188
rect 22092 19908 22148 19918
rect 22092 19814 22148 19852
rect 22540 19906 22596 19918
rect 22540 19854 22542 19906
rect 22594 19854 22596 19906
rect 21644 19294 21646 19346
rect 21698 19294 21700 19346
rect 21644 19282 21700 19294
rect 21980 19794 22036 19806
rect 21980 19742 21982 19794
rect 22034 19742 22036 19794
rect 21644 18676 21700 18686
rect 21532 18452 21588 18462
rect 21308 18340 21364 18350
rect 21308 18246 21364 18284
rect 20860 16212 20916 16828
rect 20860 16146 20916 16156
rect 20636 15262 20638 15314
rect 20690 15262 20692 15314
rect 20636 14532 20692 15262
rect 20860 15874 20916 15886
rect 20860 15822 20862 15874
rect 20914 15822 20916 15874
rect 20860 15148 20916 15822
rect 20860 15092 21028 15148
rect 20636 14476 20916 14532
rect 20524 14364 20692 14420
rect 20412 14306 20468 14318
rect 20412 14254 20414 14306
rect 20466 14254 20468 14306
rect 20412 14084 20468 14254
rect 20412 14018 20468 14028
rect 20636 13972 20692 14364
rect 20860 14308 20916 14476
rect 20860 14214 20916 14252
rect 20636 13916 20916 13972
rect 20412 13748 20468 13758
rect 20412 13074 20468 13692
rect 20748 13634 20804 13646
rect 20748 13582 20750 13634
rect 20802 13582 20804 13634
rect 20412 13022 20414 13074
rect 20466 13022 20468 13074
rect 20412 12292 20468 13022
rect 20412 12226 20468 12236
rect 20636 13300 20692 13310
rect 20524 11172 20580 11182
rect 20524 11078 20580 11116
rect 20636 9938 20692 13244
rect 20748 12962 20804 13582
rect 20748 12910 20750 12962
rect 20802 12910 20804 12962
rect 20748 12898 20804 12910
rect 20860 12068 20916 13916
rect 20972 13748 21028 15092
rect 20972 13682 21028 13692
rect 21084 13300 21140 17164
rect 21308 17780 21364 17790
rect 21308 17106 21364 17724
rect 21308 17054 21310 17106
rect 21362 17054 21364 17106
rect 21308 16996 21364 17054
rect 21532 16996 21588 18396
rect 21644 17666 21700 18620
rect 21756 18340 21812 18350
rect 21756 17778 21812 18284
rect 21756 17726 21758 17778
rect 21810 17726 21812 17778
rect 21756 17714 21812 17726
rect 21644 17614 21646 17666
rect 21698 17614 21700 17666
rect 21644 17602 21700 17614
rect 21868 17668 21924 17678
rect 21980 17668 22036 19742
rect 22540 19572 22596 19854
rect 22540 19506 22596 19516
rect 22092 19010 22148 19022
rect 22092 18958 22094 19010
rect 22146 18958 22148 19010
rect 22092 17780 22148 18958
rect 22540 19012 22596 19022
rect 22540 18918 22596 18956
rect 22988 19010 23044 19022
rect 22988 18958 22990 19010
rect 23042 18958 23044 19010
rect 22988 18788 23044 18958
rect 22988 18722 23044 18732
rect 23212 18564 23268 20132
rect 23324 20130 23380 20132
rect 23324 20078 23326 20130
rect 23378 20078 23380 20130
rect 23324 20066 23380 20078
rect 23884 19908 23940 19918
rect 23884 19906 24052 19908
rect 23884 19854 23886 19906
rect 23938 19854 24052 19906
rect 23884 19852 24052 19854
rect 23884 19842 23940 19852
rect 23324 19794 23380 19806
rect 23324 19742 23326 19794
rect 23378 19742 23380 19794
rect 23324 19234 23380 19742
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 19170 23380 19182
rect 23660 19236 23716 19246
rect 23660 19142 23716 19180
rect 23212 18498 23268 18508
rect 23548 19010 23604 19022
rect 23548 18958 23550 19010
rect 23602 18958 23604 19010
rect 23436 18340 23492 18350
rect 22092 17714 22148 17724
rect 23324 18338 23492 18340
rect 23324 18286 23438 18338
rect 23490 18286 23492 18338
rect 23324 18284 23492 18286
rect 21868 17666 22036 17668
rect 21868 17614 21870 17666
rect 21922 17614 22036 17666
rect 21868 17612 22036 17614
rect 22316 17668 22372 17678
rect 22316 17666 23156 17668
rect 22316 17614 22318 17666
rect 22370 17614 23156 17666
rect 22316 17612 23156 17614
rect 21868 17602 21924 17612
rect 22316 17602 22372 17612
rect 22988 17442 23044 17454
rect 22988 17390 22990 17442
rect 23042 17390 23044 17442
rect 21980 17220 22036 17230
rect 21756 16996 21812 17006
rect 21532 16940 21756 16996
rect 21308 16930 21364 16940
rect 21756 16902 21812 16940
rect 21980 16098 22036 17164
rect 22988 16996 23044 17390
rect 23100 17106 23156 17612
rect 23324 17220 23380 18284
rect 23436 18274 23492 18284
rect 23548 18116 23604 18958
rect 23436 18060 23604 18116
rect 23660 18564 23716 18574
rect 23436 17890 23492 18060
rect 23436 17838 23438 17890
rect 23490 17838 23492 17890
rect 23436 17826 23492 17838
rect 23548 17556 23604 17566
rect 23660 17556 23716 18508
rect 23884 18452 23940 18462
rect 23772 18450 23940 18452
rect 23772 18398 23886 18450
rect 23938 18398 23940 18450
rect 23772 18396 23940 18398
rect 23772 17668 23828 18396
rect 23884 18386 23940 18396
rect 23772 17574 23828 17612
rect 23548 17554 23716 17556
rect 23548 17502 23550 17554
rect 23602 17502 23716 17554
rect 23548 17500 23716 17502
rect 23548 17490 23604 17500
rect 23324 17164 23492 17220
rect 23100 17054 23102 17106
rect 23154 17054 23156 17106
rect 23100 17042 23156 17054
rect 21980 16046 21982 16098
rect 22034 16046 22036 16098
rect 21980 16034 22036 16046
rect 22204 16882 22260 16894
rect 22204 16830 22206 16882
rect 22258 16830 22260 16882
rect 21644 15986 21700 15998
rect 21644 15934 21646 15986
rect 21698 15934 21700 15986
rect 21644 15876 21700 15934
rect 21644 15810 21700 15820
rect 21980 15874 22036 15886
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21308 15428 21364 15438
rect 21308 15334 21364 15372
rect 21980 15428 22036 15822
rect 22204 15876 22260 16830
rect 22652 16882 22708 16894
rect 22652 16830 22654 16882
rect 22706 16830 22708 16882
rect 22428 16772 22484 16782
rect 22316 16212 22372 16222
rect 22316 16098 22372 16156
rect 22316 16046 22318 16098
rect 22370 16046 22372 16098
rect 22316 16034 22372 16046
rect 22204 15810 22260 15820
rect 21980 15362 22036 15372
rect 22428 15428 22484 16716
rect 22652 16772 22708 16830
rect 22652 16706 22708 16716
rect 22428 15362 22484 15372
rect 22988 16098 23044 16940
rect 23324 16994 23380 17006
rect 23324 16942 23326 16994
rect 23378 16942 23380 16994
rect 23324 16772 23380 16942
rect 23324 16706 23380 16716
rect 23436 16994 23492 17164
rect 23996 17108 24052 19852
rect 24220 19906 24276 19918
rect 24220 19854 24222 19906
rect 24274 19854 24276 19906
rect 24220 19796 24276 19854
rect 24668 19908 24724 19918
rect 24668 19814 24724 19852
rect 24220 19730 24276 19740
rect 24332 19124 24388 19134
rect 24108 19012 24164 19022
rect 24108 19010 24276 19012
rect 24108 18958 24110 19010
rect 24162 18958 24276 19010
rect 24108 18956 24276 18958
rect 24108 18946 24164 18956
rect 24108 18676 24164 18686
rect 24108 18582 24164 18620
rect 24220 18452 24276 18956
rect 24332 18564 24388 19068
rect 25004 19124 25060 19134
rect 25004 19030 25060 19068
rect 24332 18432 24388 18508
rect 25116 19012 25172 20132
rect 25228 19236 25284 19246
rect 25228 19142 25284 19180
rect 24444 18450 24500 18462
rect 24220 18386 24276 18396
rect 24444 18398 24446 18450
rect 24498 18398 24500 18450
rect 24444 17780 24500 18398
rect 24108 17724 24500 17780
rect 24108 17666 24164 17724
rect 24108 17614 24110 17666
rect 24162 17614 24164 17666
rect 24108 17602 24164 17614
rect 23996 17042 24052 17052
rect 24444 17106 24500 17724
rect 24780 17890 24836 17902
rect 24780 17838 24782 17890
rect 24834 17838 24836 17890
rect 24780 17668 24836 17838
rect 24780 17602 24836 17612
rect 24892 17554 24948 17566
rect 24892 17502 24894 17554
rect 24946 17502 24948 17554
rect 24444 17054 24446 17106
rect 24498 17054 24500 17106
rect 24444 17042 24500 17054
rect 24780 17442 24836 17454
rect 24780 17390 24782 17442
rect 24834 17390 24836 17442
rect 23436 16942 23438 16994
rect 23490 16942 23492 16994
rect 23212 16212 23268 16222
rect 23212 16118 23268 16156
rect 22988 16046 22990 16098
rect 23042 16046 23044 16098
rect 22988 15092 23044 16046
rect 23436 16100 23492 16942
rect 24220 16994 24276 17006
rect 24220 16942 24222 16994
rect 24274 16942 24276 16994
rect 24108 16884 24164 16894
rect 23436 16034 23492 16044
rect 23884 16882 24164 16884
rect 23884 16830 24110 16882
rect 24162 16830 24164 16882
rect 23884 16828 24164 16830
rect 23100 15988 23156 15998
rect 23100 15894 23156 15932
rect 23324 15874 23380 15886
rect 23324 15822 23326 15874
rect 23378 15822 23380 15874
rect 23324 15428 23380 15822
rect 23324 15362 23380 15372
rect 23436 15876 23492 15886
rect 23436 15202 23492 15820
rect 23884 15538 23940 16828
rect 24108 16818 24164 16828
rect 24220 16324 24276 16942
rect 24220 16258 24276 16268
rect 24668 16212 24724 16222
rect 24668 16118 24724 16156
rect 23884 15486 23886 15538
rect 23938 15486 23940 15538
rect 23884 15474 23940 15486
rect 24108 16100 24164 16110
rect 24332 16100 24388 16110
rect 24108 15538 24164 16044
rect 24108 15486 24110 15538
rect 24162 15486 24164 15538
rect 24108 15474 24164 15486
rect 24220 16044 24332 16100
rect 24220 15876 24276 16044
rect 24332 16006 24388 16044
rect 24780 16100 24836 17390
rect 24892 16882 24948 17502
rect 24892 16830 24894 16882
rect 24946 16830 24948 16882
rect 24892 16660 24948 16830
rect 24892 16594 24948 16604
rect 24780 16034 24836 16044
rect 24220 15426 24276 15820
rect 24220 15374 24222 15426
rect 24274 15374 24276 15426
rect 24220 15362 24276 15374
rect 24668 15428 24724 15438
rect 24668 15334 24724 15372
rect 25116 15428 25172 18956
rect 25116 15362 25172 15372
rect 25228 15986 25284 15998
rect 25228 15934 25230 15986
rect 25282 15934 25284 15986
rect 23436 15150 23438 15202
rect 23490 15150 23492 15202
rect 23436 15138 23492 15150
rect 22988 15026 23044 15036
rect 23548 15092 23604 15102
rect 21756 14530 21812 14542
rect 21756 14478 21758 14530
rect 21810 14478 21812 14530
rect 21420 14420 21476 14430
rect 21308 13860 21364 13870
rect 21308 13766 21364 13804
rect 21084 13234 21140 13244
rect 20860 12012 21140 12068
rect 20972 11844 21028 11854
rect 20636 9886 20638 9938
rect 20690 9886 20692 9938
rect 20524 8484 20580 8494
rect 20524 8372 20580 8428
rect 19908 7644 20356 7700
rect 20412 8370 20580 8372
rect 20412 8318 20526 8370
rect 20578 8318 20580 8370
rect 20412 8316 20580 8318
rect 19852 6804 19908 7644
rect 19404 6692 19460 6702
rect 19292 6690 19460 6692
rect 19292 6638 19406 6690
rect 19458 6638 19460 6690
rect 19292 6636 19460 6638
rect 19404 6626 19460 6636
rect 19852 6690 19908 6748
rect 19852 6638 19854 6690
rect 19906 6638 19908 6690
rect 19852 6626 19908 6638
rect 20076 6578 20132 6590
rect 20076 6526 20078 6578
rect 20130 6526 20132 6578
rect 19628 6468 19684 6478
rect 19404 6466 19684 6468
rect 19404 6414 19630 6466
rect 19682 6414 19684 6466
rect 19404 6412 19684 6414
rect 20076 6468 20132 6526
rect 20076 6412 20244 6468
rect 19404 4564 19460 6412
rect 19628 6402 19684 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19852 6132 19908 6142
rect 20188 6132 20244 6412
rect 19852 6038 19908 6076
rect 19964 6076 20244 6132
rect 19516 5124 19572 5134
rect 19516 5010 19572 5068
rect 19852 5124 19908 5134
rect 19964 5124 20020 6076
rect 20300 5796 20356 5806
rect 20412 5796 20468 8316
rect 20524 8306 20580 8316
rect 20524 7812 20580 7822
rect 20524 7140 20580 7756
rect 20636 7588 20692 9886
rect 20748 10498 20804 10510
rect 20748 10446 20750 10498
rect 20802 10446 20804 10498
rect 20748 9940 20804 10446
rect 20748 9874 20804 9884
rect 20860 10052 20916 10062
rect 20860 9938 20916 9996
rect 20860 9886 20862 9938
rect 20914 9886 20916 9938
rect 20860 9874 20916 9886
rect 20636 7522 20692 7532
rect 20748 8370 20804 8382
rect 20748 8318 20750 8370
rect 20802 8318 20804 8370
rect 20636 7364 20692 7374
rect 20636 7270 20692 7308
rect 20524 6692 20580 7084
rect 20636 6692 20692 6702
rect 20524 6690 20692 6692
rect 20524 6638 20638 6690
rect 20690 6638 20692 6690
rect 20524 6636 20692 6638
rect 20636 6626 20692 6636
rect 20748 6468 20804 8318
rect 20748 6374 20804 6412
rect 20860 8372 20916 8382
rect 20860 6244 20916 8316
rect 20972 6690 21028 11788
rect 21084 7364 21140 12012
rect 21420 10164 21476 14364
rect 21756 14308 21812 14478
rect 22428 14420 22484 14430
rect 21756 14242 21812 14252
rect 22092 14418 22484 14420
rect 22092 14366 22430 14418
rect 22482 14366 22484 14418
rect 22092 14364 22484 14366
rect 21644 14084 21700 14094
rect 21532 13860 21588 13870
rect 21532 13766 21588 13804
rect 21644 13858 21700 14028
rect 21644 13806 21646 13858
rect 21698 13806 21700 13858
rect 21644 13794 21700 13806
rect 21980 13746 22036 13758
rect 21980 13694 21982 13746
rect 22034 13694 22036 13746
rect 21980 13076 22036 13694
rect 22092 13634 22148 14364
rect 22428 14354 22484 14364
rect 22764 13860 22820 13870
rect 22092 13582 22094 13634
rect 22146 13582 22148 13634
rect 22092 13570 22148 13582
rect 22540 13858 22820 13860
rect 22540 13806 22766 13858
rect 22818 13806 22820 13858
rect 22540 13804 22820 13806
rect 21980 13010 22036 13020
rect 22316 13188 22372 13198
rect 21980 12852 22036 12862
rect 21980 12758 22036 12796
rect 22092 12738 22148 12750
rect 22092 12686 22094 12738
rect 22146 12686 22148 12738
rect 21756 12066 21812 12078
rect 21756 12014 21758 12066
rect 21810 12014 21812 12066
rect 21756 11732 21812 12014
rect 21756 11666 21812 11676
rect 22092 11620 22148 12686
rect 21868 11394 21924 11406
rect 21868 11342 21870 11394
rect 21922 11342 21924 11394
rect 21420 10108 21588 10164
rect 21196 8484 21252 8494
rect 21196 7586 21252 8428
rect 21308 8148 21364 8158
rect 21308 7698 21364 8092
rect 21420 7812 21476 10108
rect 21532 9828 21588 10108
rect 21644 10052 21700 10062
rect 21868 10052 21924 11342
rect 21700 9996 21924 10052
rect 21980 10164 22036 10174
rect 21644 9958 21700 9996
rect 21756 9828 21812 9838
rect 21532 9826 21812 9828
rect 21532 9774 21758 9826
rect 21810 9774 21812 9826
rect 21532 9772 21812 9774
rect 21756 9762 21812 9772
rect 21980 9714 22036 10108
rect 22092 9828 22148 11564
rect 22204 11172 22260 11182
rect 22204 10836 22260 11116
rect 22204 10770 22260 10780
rect 22316 10052 22372 13132
rect 22540 11618 22596 13804
rect 22764 13794 22820 13804
rect 23212 13860 23268 13870
rect 22876 13746 22932 13758
rect 22876 13694 22878 13746
rect 22930 13694 22932 13746
rect 22764 13636 22820 13646
rect 22764 13522 22820 13580
rect 22764 13470 22766 13522
rect 22818 13470 22820 13522
rect 22764 13458 22820 13470
rect 22540 11566 22542 11618
rect 22594 11566 22596 11618
rect 22540 11554 22596 11566
rect 22652 13412 22708 13422
rect 22652 12180 22708 13356
rect 22876 12964 22932 13694
rect 22988 13076 23044 13086
rect 22988 12982 23044 13020
rect 22316 9986 22372 9996
rect 22428 11170 22484 11182
rect 22428 11118 22430 11170
rect 22482 11118 22484 11170
rect 22092 9762 22148 9772
rect 22316 9828 22372 9838
rect 22316 9734 22372 9772
rect 21980 9662 21982 9714
rect 22034 9662 22036 9714
rect 21980 9650 22036 9662
rect 22428 9380 22484 11118
rect 22540 9940 22596 9950
rect 22540 9846 22596 9884
rect 22652 9828 22708 12124
rect 22764 12908 22932 12964
rect 22764 10276 22820 12908
rect 22988 12852 23044 12862
rect 22876 12738 22932 12750
rect 22876 12686 22878 12738
rect 22930 12686 22932 12738
rect 22876 11620 22932 12686
rect 22876 11060 22932 11564
rect 22876 10994 22932 11004
rect 22876 10500 22932 10510
rect 22988 10500 23044 12796
rect 23100 12740 23156 12750
rect 23212 12740 23268 13804
rect 23436 13636 23492 13646
rect 23436 12962 23492 13580
rect 23548 13634 23604 15036
rect 24444 15090 24500 15102
rect 24444 15038 24446 15090
rect 24498 15038 24500 15090
rect 24444 14756 24500 15038
rect 25116 15090 25172 15102
rect 25116 15038 25118 15090
rect 25170 15038 25172 15090
rect 24108 14700 24612 14756
rect 24108 13970 24164 14700
rect 24556 14642 24612 14700
rect 24556 14590 24558 14642
rect 24610 14590 24612 14642
rect 24556 14578 24612 14590
rect 25116 14642 25172 15038
rect 25228 15092 25284 15934
rect 25340 15148 25396 20132
rect 25564 20132 25620 20142
rect 25564 20038 25620 20076
rect 25676 20132 25844 20188
rect 25452 19010 25508 19022
rect 25452 18958 25454 19010
rect 25506 18958 25508 19010
rect 25452 17890 25508 18958
rect 25452 17838 25454 17890
rect 25506 17838 25508 17890
rect 25452 17826 25508 17838
rect 25564 19010 25620 19022
rect 25564 18958 25566 19010
rect 25618 18958 25620 19010
rect 25564 17220 25620 18958
rect 25564 17154 25620 17164
rect 25676 16996 25732 20132
rect 25900 19796 25956 22428
rect 26012 22418 26068 22428
rect 26236 23042 26292 23054
rect 26236 22990 26238 23042
rect 26290 22990 26292 23042
rect 26236 22036 26292 22990
rect 26460 22482 26516 23100
rect 26572 23044 26628 23054
rect 26572 22950 26628 22988
rect 26460 22430 26462 22482
rect 26514 22430 26516 22482
rect 26460 22418 26516 22430
rect 26236 21970 26292 21980
rect 26908 22148 26964 22158
rect 26908 21924 26964 22092
rect 26908 21858 26964 21868
rect 26348 21588 26404 21598
rect 26236 21476 26292 21486
rect 26124 21474 26292 21476
rect 26124 21422 26238 21474
rect 26290 21422 26292 21474
rect 26124 21420 26292 21422
rect 25900 19730 25956 19740
rect 26012 20020 26068 20030
rect 26012 19348 26068 19964
rect 26124 19908 26180 21420
rect 26236 21410 26292 21420
rect 26236 20804 26292 20814
rect 26236 20710 26292 20748
rect 26124 19842 26180 19852
rect 25788 19292 26068 19348
rect 25788 18116 25844 19292
rect 25900 19124 25956 19134
rect 25900 19030 25956 19068
rect 26236 19122 26292 19134
rect 26236 19070 26238 19122
rect 26290 19070 26292 19122
rect 26124 19012 26180 19022
rect 26012 19010 26180 19012
rect 26012 18958 26126 19010
rect 26178 18958 26180 19010
rect 26012 18956 26180 18958
rect 25788 18060 25956 18116
rect 25788 17892 25844 17902
rect 25788 17798 25844 17836
rect 25676 16940 25844 16996
rect 25676 16772 25732 16782
rect 25452 16770 25732 16772
rect 25452 16718 25678 16770
rect 25730 16718 25732 16770
rect 25452 16716 25732 16718
rect 25452 16100 25508 16716
rect 25676 16706 25732 16716
rect 25452 15968 25508 16044
rect 25564 15874 25620 15886
rect 25564 15822 25566 15874
rect 25618 15822 25620 15874
rect 25564 15314 25620 15822
rect 25676 15874 25732 15886
rect 25676 15822 25678 15874
rect 25730 15822 25732 15874
rect 25676 15428 25732 15822
rect 25676 15362 25732 15372
rect 25564 15262 25566 15314
rect 25618 15262 25620 15314
rect 25564 15250 25620 15262
rect 25340 15092 25508 15148
rect 25228 15026 25284 15036
rect 25116 14590 25118 14642
rect 25170 14590 25172 14642
rect 25116 14578 25172 14590
rect 25228 14420 25284 14430
rect 24108 13918 24110 13970
rect 24162 13918 24164 13970
rect 24108 13906 24164 13918
rect 24220 14308 24276 14318
rect 25228 14308 25284 14364
rect 23548 13582 23550 13634
rect 23602 13582 23604 13634
rect 23548 13412 23604 13582
rect 23548 13346 23604 13356
rect 23660 13524 23716 13534
rect 23436 12910 23438 12962
rect 23490 12910 23492 12962
rect 23436 12898 23492 12910
rect 23100 12738 23268 12740
rect 23100 12686 23102 12738
rect 23154 12686 23268 12738
rect 23100 12684 23268 12686
rect 23100 12674 23156 12684
rect 23212 11508 23268 12684
rect 23660 12180 23716 13468
rect 23660 12048 23716 12124
rect 24220 12962 24276 14252
rect 25116 14306 25284 14308
rect 25116 14254 25230 14306
rect 25282 14254 25284 14306
rect 25116 14252 25284 14254
rect 24780 13858 24836 13870
rect 24780 13806 24782 13858
rect 24834 13806 24836 13858
rect 24220 12910 24222 12962
rect 24274 12910 24276 12962
rect 22876 10498 23156 10500
rect 22876 10446 22878 10498
rect 22930 10446 23156 10498
rect 22876 10444 23156 10446
rect 22876 10434 22932 10444
rect 22764 10210 22820 10220
rect 22652 9826 22932 9828
rect 22652 9774 22654 9826
rect 22706 9774 22932 9826
rect 22652 9772 22932 9774
rect 22652 9762 22708 9772
rect 22876 9492 22932 9772
rect 22428 9314 22484 9324
rect 22764 9436 22932 9492
rect 22988 9492 23044 9502
rect 22316 9156 22372 9166
rect 21644 8932 21700 8942
rect 21644 8148 21700 8876
rect 21756 8930 21812 8942
rect 21756 8878 21758 8930
rect 21810 8878 21812 8930
rect 21756 8372 21812 8878
rect 22092 8372 22148 8382
rect 21756 8370 22148 8372
rect 21756 8318 22094 8370
rect 22146 8318 22148 8370
rect 21756 8316 22148 8318
rect 22092 8306 22148 8316
rect 22316 8258 22372 9100
rect 22428 9042 22484 9054
rect 22428 8990 22430 9042
rect 22482 8990 22484 9042
rect 22428 8372 22484 8990
rect 22428 8306 22484 8316
rect 22540 9044 22596 9054
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8194 22372 8206
rect 21756 8148 21812 8158
rect 22204 8148 22260 8158
rect 21420 7746 21476 7756
rect 21532 8146 21812 8148
rect 21532 8094 21758 8146
rect 21810 8094 21812 8146
rect 21532 8092 21812 8094
rect 21308 7646 21310 7698
rect 21362 7646 21364 7698
rect 21308 7634 21364 7646
rect 21196 7534 21198 7586
rect 21250 7534 21252 7586
rect 21196 7522 21252 7534
rect 21420 7586 21476 7598
rect 21420 7534 21422 7586
rect 21474 7534 21476 7586
rect 21420 7476 21476 7534
rect 21308 7420 21476 7476
rect 21308 7364 21364 7420
rect 21084 7308 21308 7364
rect 20972 6638 20974 6690
rect 21026 6638 21028 6690
rect 20972 6626 21028 6638
rect 20300 5794 20468 5796
rect 20300 5742 20302 5794
rect 20354 5742 20468 5794
rect 20300 5740 20468 5742
rect 20748 6188 20916 6244
rect 20300 5730 20356 5740
rect 19852 5122 20020 5124
rect 19852 5070 19854 5122
rect 19906 5070 20020 5122
rect 19852 5068 20020 5070
rect 20300 5348 20356 5358
rect 19852 5058 19908 5068
rect 19516 4958 19518 5010
rect 19570 4958 19572 5010
rect 19516 4946 19572 4958
rect 19628 5012 19684 5022
rect 19628 4918 19684 4956
rect 20300 5010 20356 5292
rect 20300 4958 20302 5010
rect 20354 4958 20356 5010
rect 20300 4946 20356 4958
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19404 4508 20020 4564
rect 19964 4450 20020 4508
rect 19964 4398 19966 4450
rect 20018 4398 20020 4450
rect 19964 4386 20020 4398
rect 20748 4338 20804 6188
rect 20860 5236 20916 5246
rect 20860 5142 20916 5180
rect 20748 4286 20750 4338
rect 20802 4286 20804 4338
rect 20748 4274 20804 4286
rect 21308 4228 21364 7308
rect 21308 4162 21364 4172
rect 21420 6804 21476 6814
rect 21308 4004 21364 4014
rect 20188 3666 20244 3678
rect 20188 3614 20190 3666
rect 20242 3614 20244 3666
rect 19404 3556 19460 3566
rect 19180 3554 19460 3556
rect 19180 3502 19406 3554
rect 19458 3502 19460 3554
rect 19180 3500 19460 3502
rect 19404 3490 19460 3500
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 2996 20244 3614
rect 19964 2940 20244 2996
rect 19964 800 20020 2940
rect 21308 800 21364 3948
rect 21420 3778 21476 6748
rect 21532 6692 21588 8092
rect 21756 8082 21812 8092
rect 22092 8146 22260 8148
rect 22092 8094 22206 8146
rect 22258 8094 22260 8146
rect 22092 8092 22260 8094
rect 21980 8034 22036 8046
rect 21980 7982 21982 8034
rect 22034 7982 22036 8034
rect 21532 5236 21588 6636
rect 21756 7924 21812 7934
rect 21532 5170 21588 5180
rect 21644 6578 21700 6590
rect 21644 6526 21646 6578
rect 21698 6526 21700 6578
rect 21644 5124 21700 6526
rect 21644 5058 21700 5068
rect 21756 5122 21812 7868
rect 21980 7812 22036 7982
rect 22092 8036 22148 8092
rect 22204 8082 22260 8092
rect 22092 7970 22148 7980
rect 22036 7756 22148 7812
rect 21980 7746 22036 7756
rect 22092 7586 22148 7756
rect 22092 7534 22094 7586
rect 22146 7534 22148 7586
rect 22092 7522 22148 7534
rect 22428 7588 22484 7598
rect 22540 7588 22596 8988
rect 22428 7586 22596 7588
rect 22428 7534 22430 7586
rect 22482 7534 22596 7586
rect 22428 7532 22596 7534
rect 22428 7522 22484 7532
rect 22764 7252 22820 9436
rect 22988 9044 23044 9436
rect 22988 8950 23044 8988
rect 23100 8932 23156 10444
rect 23212 9828 23268 11452
rect 23548 11844 23604 11854
rect 23548 10834 23604 11788
rect 23548 10782 23550 10834
rect 23602 10782 23604 10834
rect 23548 10770 23604 10782
rect 23884 11732 23940 11742
rect 23436 10724 23492 10734
rect 23436 10630 23492 10668
rect 23212 9762 23268 9772
rect 23660 10388 23716 10398
rect 23436 9604 23492 9614
rect 23100 8866 23156 8876
rect 23324 9602 23492 9604
rect 23324 9550 23438 9602
rect 23490 9550 23492 9602
rect 23324 9548 23492 9550
rect 22652 7196 22820 7252
rect 22876 8372 22932 8382
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5058 21812 5070
rect 22204 6580 22260 6590
rect 22204 5796 22260 6524
rect 22428 6468 22484 6478
rect 22428 6018 22484 6412
rect 22652 6132 22708 7196
rect 22764 6692 22820 6702
rect 22764 6598 22820 6636
rect 22652 6066 22708 6076
rect 22428 5966 22430 6018
rect 22482 5966 22484 6018
rect 22428 5954 22484 5966
rect 22876 5908 22932 8316
rect 23100 8036 23156 8046
rect 23100 7698 23156 7980
rect 23100 7646 23102 7698
rect 23154 7646 23156 7698
rect 23100 7634 23156 7646
rect 22988 7474 23044 7486
rect 22988 7422 22990 7474
rect 23042 7422 23044 7474
rect 22988 6692 23044 7422
rect 23212 7362 23268 7374
rect 23212 7310 23214 7362
rect 23266 7310 23268 7362
rect 23212 7140 23268 7310
rect 23212 7074 23268 7084
rect 22988 6626 23044 6636
rect 23212 6692 23268 6702
rect 23324 6692 23380 9548
rect 23436 9538 23492 9548
rect 23548 9602 23604 9614
rect 23548 9550 23550 9602
rect 23602 9550 23604 9602
rect 23548 9268 23604 9550
rect 23660 9492 23716 10332
rect 23772 9828 23828 9838
rect 23772 9734 23828 9772
rect 23660 9436 23828 9492
rect 23548 9202 23604 9212
rect 23436 9042 23492 9054
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23436 8820 23492 8990
rect 23548 9044 23604 9054
rect 23548 8950 23604 8988
rect 23660 9042 23716 9054
rect 23660 8990 23662 9042
rect 23714 8990 23716 9042
rect 23660 8932 23716 8990
rect 23660 8866 23716 8876
rect 23436 8764 23604 8820
rect 23548 8484 23604 8764
rect 23548 7476 23604 8428
rect 23772 7588 23828 9436
rect 23884 8258 23940 11676
rect 24220 11506 24276 12910
rect 24444 13748 24500 13758
rect 24220 11454 24222 11506
rect 24274 11454 24276 11506
rect 24220 11442 24276 11454
rect 24332 12740 24388 12750
rect 24332 11844 24388 12684
rect 24332 10834 24388 11788
rect 24332 10782 24334 10834
rect 24386 10782 24388 10834
rect 24332 10770 24388 10782
rect 24220 10610 24276 10622
rect 24220 10558 24222 10610
rect 24274 10558 24276 10610
rect 23996 9716 24052 9726
rect 23996 9622 24052 9660
rect 23884 8206 23886 8258
rect 23938 8206 23940 8258
rect 23884 8194 23940 8206
rect 23996 9380 24052 9390
rect 23884 7588 23940 7598
rect 23772 7586 23940 7588
rect 23772 7534 23886 7586
rect 23938 7534 23940 7586
rect 23772 7532 23940 7534
rect 23884 7522 23940 7532
rect 23660 7476 23716 7486
rect 23548 7420 23660 7476
rect 23660 7382 23716 7420
rect 23436 7250 23492 7262
rect 23436 7198 23438 7250
rect 23490 7198 23492 7250
rect 23436 6916 23492 7198
rect 23996 6916 24052 9324
rect 24108 9044 24164 9054
rect 24108 8950 24164 8988
rect 24220 8820 24276 10558
rect 24444 10388 24500 13692
rect 24780 13748 24836 13806
rect 24780 13682 24836 13692
rect 24892 13746 24948 13758
rect 24892 13694 24894 13746
rect 24946 13694 24948 13746
rect 24556 13636 24612 13646
rect 24556 10722 24612 13580
rect 24780 13522 24836 13534
rect 24780 13470 24782 13522
rect 24834 13470 24836 13522
rect 24668 13412 24724 13422
rect 24668 10836 24724 13356
rect 24668 10770 24724 10780
rect 24556 10670 24558 10722
rect 24610 10670 24612 10722
rect 24556 10658 24612 10670
rect 24780 10610 24836 13470
rect 24892 13412 24948 13694
rect 24892 12852 24948 13356
rect 24892 12786 24948 12796
rect 25004 12850 25060 12862
rect 25004 12798 25006 12850
rect 25058 12798 25060 12850
rect 24780 10558 24782 10610
rect 24834 10558 24836 10610
rect 24780 10546 24836 10558
rect 24668 10498 24724 10510
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10388 24724 10446
rect 25004 10388 25060 12798
rect 24668 10332 25060 10388
rect 24444 10322 24500 10332
rect 25004 10164 25060 10174
rect 24668 9938 24724 9950
rect 24668 9886 24670 9938
rect 24722 9886 24724 9938
rect 24556 9714 24612 9726
rect 24556 9662 24558 9714
rect 24610 9662 24612 9714
rect 24556 9380 24612 9662
rect 24556 9266 24612 9324
rect 24556 9214 24558 9266
rect 24610 9214 24612 9266
rect 24556 9202 24612 9214
rect 24668 9156 24724 9886
rect 25004 9714 25060 10108
rect 25004 9662 25006 9714
rect 25058 9662 25060 9714
rect 25004 9650 25060 9662
rect 24780 9602 24836 9614
rect 24780 9550 24782 9602
rect 24834 9550 24836 9602
rect 24780 9492 24836 9550
rect 25116 9492 25172 14252
rect 25228 14242 25284 14252
rect 25452 13972 25508 15092
rect 25452 13748 25508 13916
rect 24780 9436 25172 9492
rect 25340 12180 25396 12190
rect 24668 9090 24724 9100
rect 24780 9044 24836 9054
rect 24780 8950 24836 8988
rect 24220 8754 24276 8764
rect 24668 8930 24724 8942
rect 24668 8878 24670 8930
rect 24722 8878 24724 8930
rect 24668 8820 24724 8878
rect 24668 8754 24724 8764
rect 24332 8708 24388 8718
rect 24108 6916 24164 6926
rect 23436 6860 23604 6916
rect 23996 6914 24164 6916
rect 23996 6862 24110 6914
rect 24162 6862 24164 6914
rect 23996 6860 24164 6862
rect 23548 6804 23604 6860
rect 24108 6850 24164 6860
rect 23548 6748 23828 6804
rect 23212 6690 23380 6692
rect 23212 6638 23214 6690
rect 23266 6638 23380 6690
rect 23212 6636 23380 6638
rect 23436 6692 23492 6702
rect 23436 6690 23716 6692
rect 23436 6638 23438 6690
rect 23490 6638 23716 6690
rect 23436 6636 23716 6638
rect 23212 6626 23268 6636
rect 23436 6626 23492 6636
rect 22988 6466 23044 6478
rect 22988 6414 22990 6466
rect 23042 6414 23044 6466
rect 22988 6356 23044 6414
rect 23100 6468 23156 6478
rect 23100 6374 23156 6412
rect 23436 6468 23492 6478
rect 22988 6290 23044 6300
rect 23100 5908 23156 5918
rect 22876 5906 23156 5908
rect 22876 5854 23102 5906
rect 23154 5854 23156 5906
rect 22876 5852 23156 5854
rect 22204 4228 22260 5740
rect 22204 4162 22260 4172
rect 22316 5234 22372 5246
rect 22316 5182 22318 5234
rect 22370 5182 22372 5234
rect 22316 4004 22372 5182
rect 23100 4900 23156 5852
rect 23100 4834 23156 4844
rect 23436 4450 23492 6412
rect 23660 6130 23716 6636
rect 23772 6244 23828 6748
rect 24108 6692 24164 6702
rect 23996 6580 24052 6590
rect 23772 6178 23828 6188
rect 23884 6578 24052 6580
rect 23884 6526 23998 6578
rect 24050 6526 24052 6578
rect 23884 6524 24052 6526
rect 23660 6078 23662 6130
rect 23714 6078 23716 6130
rect 23660 6066 23716 6078
rect 23772 5908 23828 5918
rect 23548 5906 23828 5908
rect 23548 5854 23774 5906
rect 23826 5854 23828 5906
rect 23548 5852 23828 5854
rect 23548 5012 23604 5852
rect 23772 5842 23828 5852
rect 23660 5684 23716 5694
rect 23660 5346 23716 5628
rect 23884 5348 23940 6524
rect 23996 6514 24052 6524
rect 23996 6020 24052 6030
rect 23996 5906 24052 5964
rect 23996 5854 23998 5906
rect 24050 5854 24052 5906
rect 23996 5842 24052 5854
rect 24108 5460 24164 6636
rect 24220 6468 24276 6478
rect 24332 6468 24388 8652
rect 24668 8596 24724 8606
rect 24444 7364 24500 7374
rect 24444 7270 24500 7308
rect 24668 7362 24724 8540
rect 25228 8372 25284 8382
rect 25228 8278 25284 8316
rect 25340 7700 25396 12124
rect 25452 11508 25508 13692
rect 25564 14868 25620 14878
rect 25564 12404 25620 14812
rect 25788 13972 25844 16940
rect 25900 16884 25956 18060
rect 26012 17780 26068 18956
rect 26124 18946 26180 18956
rect 26124 18452 26180 18462
rect 26124 18358 26180 18396
rect 26236 17892 26292 19070
rect 26236 17826 26292 17836
rect 26012 17686 26068 17724
rect 26236 17444 26292 17454
rect 26236 17106 26292 17388
rect 26348 17220 26404 21532
rect 26684 21588 26740 21598
rect 26684 21494 26740 21532
rect 26572 20692 26628 20702
rect 26572 20598 26628 20636
rect 27020 20580 27076 24556
rect 28028 24052 28084 24062
rect 28028 23958 28084 23996
rect 30044 23940 30100 27020
rect 36316 27076 36372 27086
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 33068 25284 33124 25294
rect 30492 24724 30548 24734
rect 30156 24612 30212 24622
rect 30156 24610 30324 24612
rect 30156 24558 30158 24610
rect 30210 24558 30324 24610
rect 30156 24556 30324 24558
rect 30156 24546 30212 24556
rect 30044 23884 30212 23940
rect 28700 23714 28756 23726
rect 28700 23662 28702 23714
rect 28754 23662 28756 23714
rect 28700 23268 28756 23662
rect 28700 23202 28756 23212
rect 29596 23714 29652 23726
rect 29596 23662 29598 23714
rect 29650 23662 29652 23714
rect 27132 23042 27188 23054
rect 27132 22990 27134 23042
rect 27186 22990 27188 23042
rect 27132 21700 27188 22990
rect 27580 23044 27636 23054
rect 28252 23044 28308 23054
rect 27580 23042 27972 23044
rect 27580 22990 27582 23042
rect 27634 22990 27972 23042
rect 27580 22988 27972 22990
rect 27580 22978 27636 22988
rect 27804 22260 27860 22270
rect 27804 22166 27860 22204
rect 27468 22148 27524 22158
rect 27468 22146 27748 22148
rect 27468 22094 27470 22146
rect 27522 22094 27748 22146
rect 27468 22092 27748 22094
rect 27468 22082 27524 22092
rect 27132 21634 27188 21644
rect 27020 20486 27076 20524
rect 27132 21474 27188 21486
rect 27580 21476 27636 21486
rect 27132 21422 27134 21474
rect 27186 21422 27188 21474
rect 27132 20132 27188 21422
rect 27132 20066 27188 20076
rect 27356 21474 27636 21476
rect 27356 21422 27582 21474
rect 27634 21422 27636 21474
rect 27356 21420 27636 21422
rect 26572 19906 26628 19918
rect 26572 19854 26574 19906
rect 26626 19854 26628 19906
rect 26572 18676 26628 19854
rect 26908 19906 26964 19918
rect 26908 19854 26910 19906
rect 26962 19854 26964 19906
rect 26908 19796 26964 19854
rect 26908 19730 26964 19740
rect 27356 19684 27412 21420
rect 27580 21410 27636 21420
rect 27580 20580 27636 20590
rect 27356 19618 27412 19628
rect 27468 19906 27524 19918
rect 27468 19854 27470 19906
rect 27522 19854 27524 19906
rect 27132 19460 27188 19470
rect 26572 18610 26628 18620
rect 26684 19010 26740 19022
rect 26684 18958 26686 19010
rect 26738 18958 26740 19010
rect 26684 18452 26740 18958
rect 27132 19012 27188 19404
rect 27468 19348 27524 19854
rect 27132 18918 27188 18956
rect 27244 19292 27524 19348
rect 27132 18676 27188 18686
rect 26684 18386 26740 18396
rect 27020 18452 27076 18462
rect 26796 18338 26852 18350
rect 26796 18286 26798 18338
rect 26850 18286 26852 18338
rect 26572 17556 26628 17566
rect 26572 17462 26628 17500
rect 26684 17444 26740 17454
rect 26684 17350 26740 17388
rect 26348 17164 26740 17220
rect 26236 17054 26238 17106
rect 26290 17054 26292 17106
rect 26236 17042 26292 17054
rect 26460 16996 26516 17006
rect 25900 16828 26292 16884
rect 25900 16660 25956 16670
rect 25900 16100 25956 16604
rect 25900 16006 25956 16044
rect 26012 15986 26068 15998
rect 26012 15934 26014 15986
rect 26066 15934 26068 15986
rect 25900 15540 25956 15550
rect 26012 15540 26068 15934
rect 26236 15988 26292 16828
rect 26348 16212 26404 16222
rect 26348 16118 26404 16156
rect 26236 15932 26404 15988
rect 25900 15538 26068 15540
rect 25900 15486 25902 15538
rect 25954 15486 26068 15538
rect 25900 15484 26068 15486
rect 26236 15764 26292 15774
rect 25900 15474 25956 15484
rect 26236 15426 26292 15708
rect 26236 15374 26238 15426
rect 26290 15374 26292 15426
rect 26236 15362 26292 15374
rect 26012 15316 26068 15326
rect 26012 15222 26068 15260
rect 26348 14868 26404 15932
rect 26348 14802 26404 14812
rect 25900 14532 25956 14542
rect 25900 14308 25956 14476
rect 26460 14418 26516 16940
rect 26572 16884 26628 16894
rect 26572 14532 26628 16828
rect 26572 14466 26628 14476
rect 26460 14366 26462 14418
rect 26514 14366 26516 14418
rect 26460 14354 26516 14366
rect 25900 14214 25956 14252
rect 26572 14306 26628 14318
rect 26572 14254 26574 14306
rect 26626 14254 26628 14306
rect 25788 13916 26068 13972
rect 25676 13748 25732 13758
rect 25676 13654 25732 13692
rect 25900 13748 25956 13758
rect 25900 13654 25956 13692
rect 25788 13636 25844 13646
rect 25788 13542 25844 13580
rect 26012 13300 26068 13916
rect 26348 13748 26404 13758
rect 26348 13654 26404 13692
rect 26236 13300 26292 13310
rect 26012 13244 26236 13300
rect 26012 13076 26068 13086
rect 25900 12740 25956 12750
rect 25564 12348 25732 12404
rect 25452 11442 25508 11452
rect 25564 12178 25620 12190
rect 25564 12126 25566 12178
rect 25618 12126 25620 12178
rect 25452 10388 25508 10398
rect 25452 9938 25508 10332
rect 25564 10164 25620 12126
rect 25676 10610 25732 12348
rect 25788 12290 25844 12302
rect 25788 12238 25790 12290
rect 25842 12238 25844 12290
rect 25788 11396 25844 12238
rect 25900 12290 25956 12684
rect 25900 12238 25902 12290
rect 25954 12238 25956 12290
rect 25900 12226 25956 12238
rect 25788 11330 25844 11340
rect 25900 11508 25956 11518
rect 25900 11172 25956 11452
rect 25676 10558 25678 10610
rect 25730 10558 25732 10610
rect 25676 10500 25732 10558
rect 25676 10434 25732 10444
rect 25788 11116 25956 11172
rect 25564 10098 25620 10108
rect 25452 9886 25454 9938
rect 25506 9886 25508 9938
rect 25452 9874 25508 9886
rect 25676 10052 25732 10062
rect 25564 9716 25620 9726
rect 25564 9266 25620 9660
rect 25564 9214 25566 9266
rect 25618 9214 25620 9266
rect 25564 9202 25620 9214
rect 25676 9380 25732 9996
rect 25676 9266 25732 9324
rect 25676 9214 25678 9266
rect 25730 9214 25732 9266
rect 25676 9202 25732 9214
rect 25676 8932 25732 8942
rect 25564 7700 25620 7710
rect 25340 7698 25620 7700
rect 25340 7646 25566 7698
rect 25618 7646 25620 7698
rect 25340 7644 25620 7646
rect 25564 7634 25620 7644
rect 24668 7310 24670 7362
rect 24722 7310 24724 7362
rect 24668 6804 24724 7310
rect 24668 6738 24724 6748
rect 24780 7588 24836 7598
rect 24668 6580 24724 6590
rect 24556 6578 24724 6580
rect 24556 6526 24670 6578
rect 24722 6526 24724 6578
rect 24556 6524 24724 6526
rect 24220 6466 24388 6468
rect 24220 6414 24222 6466
rect 24274 6414 24388 6466
rect 24220 6412 24388 6414
rect 24220 6402 24276 6412
rect 24220 6244 24276 6254
rect 24220 5682 24276 6188
rect 24220 5630 24222 5682
rect 24274 5630 24276 5682
rect 24220 5572 24276 5630
rect 24220 5506 24276 5516
rect 23660 5294 23662 5346
rect 23714 5294 23716 5346
rect 23660 5282 23716 5294
rect 23772 5292 23940 5348
rect 23996 5404 24164 5460
rect 23548 4946 23604 4956
rect 23772 4898 23828 5292
rect 23996 5236 24052 5404
rect 24220 5348 24276 5358
rect 24220 5254 24276 5292
rect 23884 5124 23940 5134
rect 23996 5124 24052 5180
rect 23884 5122 24052 5124
rect 23884 5070 23886 5122
rect 23938 5070 24052 5122
rect 23884 5068 24052 5070
rect 24108 5124 24164 5134
rect 24108 5122 24276 5124
rect 24108 5070 24110 5122
rect 24162 5070 24276 5122
rect 24108 5068 24276 5070
rect 23884 5058 23940 5068
rect 24108 5058 24164 5068
rect 24220 5012 24276 5068
rect 23772 4846 23774 4898
rect 23826 4846 23828 4898
rect 23772 4834 23828 4846
rect 24108 4900 24164 4910
rect 23436 4398 23438 4450
rect 23490 4398 23492 4450
rect 23436 4386 23492 4398
rect 23996 4788 24052 4798
rect 22316 3938 22372 3948
rect 21420 3726 21422 3778
rect 21474 3726 21476 3778
rect 21420 3714 21476 3726
rect 23996 3780 24052 4732
rect 24108 4340 24164 4844
rect 24108 4208 24164 4284
rect 21532 3668 21588 3678
rect 21532 3574 21588 3612
rect 22540 3444 22596 3454
rect 22540 3442 22708 3444
rect 22540 3390 22542 3442
rect 22594 3390 22708 3442
rect 22540 3388 22708 3390
rect 22540 3378 22596 3388
rect 22652 2996 22708 3388
rect 22652 800 22708 2940
rect 23996 800 24052 3724
rect 24220 3668 24276 4956
rect 24220 3602 24276 3612
rect 24332 3666 24388 6412
rect 24444 6466 24500 6478
rect 24444 6414 24446 6466
rect 24498 6414 24500 6466
rect 24444 6132 24500 6414
rect 24444 6066 24500 6076
rect 24444 5908 24500 5918
rect 24444 5814 24500 5852
rect 24332 3614 24334 3666
rect 24386 3614 24388 3666
rect 24332 3602 24388 3614
rect 24556 3388 24612 6524
rect 24668 6514 24724 6524
rect 24780 5906 24836 7532
rect 24780 5854 24782 5906
rect 24834 5854 24836 5906
rect 24780 5842 24836 5854
rect 24892 7364 24948 7374
rect 24892 7028 24948 7308
rect 24892 5908 24948 6972
rect 24892 5842 24948 5852
rect 25004 6804 25060 6814
rect 25004 5346 25060 6748
rect 25452 6692 25508 6702
rect 25452 6598 25508 6636
rect 25676 6690 25732 8876
rect 25788 8708 25844 11116
rect 25900 10724 25956 10734
rect 26012 10724 26068 13020
rect 25956 10668 26068 10724
rect 26124 10836 26180 10846
rect 25900 10630 25956 10668
rect 25900 10500 25956 10510
rect 25900 9266 25956 10444
rect 26012 10388 26068 10398
rect 26124 10388 26180 10780
rect 26068 10332 26180 10388
rect 26012 9826 26068 10332
rect 26012 9774 26014 9826
rect 26066 9774 26068 9826
rect 26012 9762 26068 9774
rect 25900 9214 25902 9266
rect 25954 9214 25956 9266
rect 25900 9202 25956 9214
rect 25788 8642 25844 8652
rect 26124 9156 26180 9166
rect 26124 8260 26180 9100
rect 26124 8194 26180 8204
rect 26236 8820 26292 13244
rect 26572 12852 26628 14254
rect 26572 12786 26628 12796
rect 26684 12628 26740 17164
rect 26796 16322 26852 18286
rect 26908 17556 26964 17566
rect 26908 17462 26964 17500
rect 27020 16884 27076 18396
rect 27020 16752 27076 16828
rect 26796 16270 26798 16322
rect 26850 16270 26852 16322
rect 26796 16258 26852 16270
rect 27020 16100 27076 16110
rect 27132 16100 27188 18620
rect 27244 17332 27300 19292
rect 27356 17892 27412 17902
rect 27356 17798 27412 17836
rect 27468 17556 27524 17566
rect 27468 17462 27524 17500
rect 27244 16996 27300 17276
rect 27244 16930 27300 16940
rect 27468 16548 27524 16558
rect 27356 16436 27412 16446
rect 27356 16210 27412 16380
rect 27356 16158 27358 16210
rect 27410 16158 27412 16210
rect 27356 16146 27412 16158
rect 27020 16098 27188 16100
rect 27020 16046 27022 16098
rect 27074 16046 27188 16098
rect 27020 16044 27188 16046
rect 27244 16098 27300 16110
rect 27244 16046 27246 16098
rect 27298 16046 27300 16098
rect 27020 15764 27076 16044
rect 27020 15698 27076 15708
rect 26908 15652 26964 15662
rect 26908 15538 26964 15596
rect 26908 15486 26910 15538
rect 26962 15486 26964 15538
rect 26908 15474 26964 15486
rect 27132 15540 27188 15550
rect 27132 15446 27188 15484
rect 26796 15316 26852 15326
rect 26796 15222 26852 15260
rect 27244 15204 27300 16046
rect 27468 16098 27524 16492
rect 27468 16046 27470 16098
rect 27522 16046 27524 16098
rect 27468 16034 27524 16046
rect 27244 15138 27300 15148
rect 27356 15988 27412 15998
rect 27020 15092 27076 15102
rect 27020 13970 27076 15036
rect 27244 14756 27300 14766
rect 27356 14756 27412 15932
rect 27468 15316 27524 15326
rect 27468 15222 27524 15260
rect 27244 14754 27412 14756
rect 27244 14702 27246 14754
rect 27298 14702 27412 14754
rect 27244 14700 27412 14702
rect 27244 14690 27300 14700
rect 27132 14532 27188 14542
rect 27188 14476 27412 14532
rect 27132 14438 27188 14476
rect 27244 14308 27300 14318
rect 27244 14214 27300 14252
rect 27020 13918 27022 13970
rect 27074 13918 27076 13970
rect 27020 13906 27076 13918
rect 27244 13972 27300 13982
rect 26796 13746 26852 13758
rect 26796 13694 26798 13746
rect 26850 13694 26852 13746
rect 26796 13076 26852 13694
rect 26908 13748 26964 13758
rect 26908 13654 26964 13692
rect 26796 13010 26852 13020
rect 27132 13076 27188 13086
rect 27132 12982 27188 13020
rect 26684 12562 26740 12572
rect 26908 12180 26964 12190
rect 27244 12180 27300 13916
rect 27356 13748 27412 14476
rect 27356 13616 27412 13692
rect 27580 13524 27636 20524
rect 27692 19684 27748 22092
rect 27916 21252 27972 22988
rect 28140 23042 28308 23044
rect 28140 22990 28254 23042
rect 28306 22990 28308 23042
rect 28140 22988 28308 22990
rect 28028 21476 28084 21486
rect 28028 21382 28084 21420
rect 27916 21196 28084 21252
rect 27804 21028 27860 21038
rect 27804 20188 27860 20972
rect 27916 20578 27972 20590
rect 27916 20526 27918 20578
rect 27970 20526 27972 20578
rect 27916 20468 27972 20526
rect 27916 20402 27972 20412
rect 27804 20132 27972 20188
rect 27804 20020 27860 20030
rect 27804 19926 27860 19964
rect 27692 19618 27748 19628
rect 27916 19460 27972 20132
rect 27692 19404 27972 19460
rect 27692 19346 27748 19404
rect 27692 19294 27694 19346
rect 27746 19294 27748 19346
rect 27692 19282 27748 19294
rect 27916 17220 27972 19404
rect 28028 19460 28084 21196
rect 28140 21028 28196 22988
rect 28252 22978 28308 22988
rect 28588 23042 28644 23054
rect 28588 22990 28590 23042
rect 28642 22990 28644 23042
rect 28588 22932 28644 22990
rect 28588 22866 28644 22876
rect 29372 23042 29428 23054
rect 29372 22990 29374 23042
rect 29426 22990 29428 23042
rect 28140 20962 28196 20972
rect 28252 22596 28308 22606
rect 28252 20188 28308 22540
rect 28812 22484 28868 22494
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28476 21474 28532 21486
rect 28476 21422 28478 21474
rect 28530 21422 28532 21474
rect 28364 20578 28420 20590
rect 28364 20526 28366 20578
rect 28418 20526 28420 20578
rect 28364 20356 28420 20526
rect 28364 20290 28420 20300
rect 28252 20132 28420 20188
rect 28028 19394 28084 19404
rect 28140 20020 28196 20030
rect 28140 19908 28196 19964
rect 28252 19908 28308 19918
rect 28140 19906 28308 19908
rect 28140 19854 28254 19906
rect 28306 19854 28308 19906
rect 28140 19852 28308 19854
rect 28140 19348 28196 19852
rect 28252 19842 28308 19852
rect 28140 19282 28196 19292
rect 28252 19684 28308 19694
rect 28028 19236 28084 19246
rect 28028 17892 28084 19180
rect 28140 19010 28196 19022
rect 28140 18958 28142 19010
rect 28194 18958 28196 19010
rect 28140 18564 28196 18958
rect 28140 18498 28196 18508
rect 28140 17892 28196 17902
rect 28028 17890 28196 17892
rect 28028 17838 28142 17890
rect 28194 17838 28196 17890
rect 28028 17836 28196 17838
rect 28028 17554 28084 17566
rect 28028 17502 28030 17554
rect 28082 17502 28084 17554
rect 28028 17444 28084 17502
rect 28028 17378 28084 17388
rect 27916 17164 28084 17220
rect 27804 16770 27860 16782
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27804 16436 27860 16718
rect 27804 16370 27860 16380
rect 28028 16098 28084 17164
rect 28028 16046 28030 16098
rect 28082 16046 28084 16098
rect 28028 15092 28084 16046
rect 28140 15540 28196 17836
rect 28252 16436 28308 19628
rect 28364 16884 28420 20132
rect 28476 16996 28532 21422
rect 28588 20580 28644 22094
rect 28812 21812 28868 22428
rect 29372 21924 29428 22990
rect 29484 22484 29540 22494
rect 29484 22390 29540 22428
rect 29372 21858 29428 21868
rect 28812 21680 28868 21756
rect 29260 21474 29316 21486
rect 29260 21422 29262 21474
rect 29314 21422 29316 21474
rect 28700 20692 28756 20702
rect 28700 20598 28756 20636
rect 28588 20514 28644 20524
rect 29260 20188 29316 21422
rect 29596 20916 29652 23662
rect 30044 23714 30100 23726
rect 30044 23662 30046 23714
rect 30098 23662 30100 23714
rect 29708 23156 29764 23166
rect 29708 23062 29764 23100
rect 30044 22932 30100 23662
rect 30044 22866 30100 22876
rect 29596 20850 29652 20860
rect 29932 22708 29988 22718
rect 29932 20914 29988 22652
rect 30044 22484 30100 22494
rect 30156 22484 30212 23884
rect 30044 22482 30212 22484
rect 30044 22430 30046 22482
rect 30098 22430 30212 22482
rect 30044 22428 30212 22430
rect 30044 22372 30100 22428
rect 30044 22306 30100 22316
rect 30268 22260 30324 24556
rect 30492 24050 30548 24668
rect 30604 24612 30660 24622
rect 30604 24518 30660 24556
rect 31836 24610 31892 24622
rect 31836 24558 31838 24610
rect 31890 24558 31892 24610
rect 30492 23998 30494 24050
rect 30546 23998 30548 24050
rect 30492 23604 30548 23998
rect 31164 23714 31220 23726
rect 31164 23662 31166 23714
rect 31218 23662 31220 23714
rect 31164 23548 31220 23662
rect 30492 23538 30548 23548
rect 30828 23492 31220 23548
rect 31500 23714 31556 23726
rect 31500 23662 31502 23714
rect 31554 23662 31556 23714
rect 30828 23156 30884 23492
rect 30492 23042 30548 23054
rect 30492 22990 30494 23042
rect 30546 22990 30548 23042
rect 30492 22596 30548 22990
rect 30828 23042 30884 23100
rect 30828 22990 30830 23042
rect 30882 22990 30884 23042
rect 30492 22530 30548 22540
rect 30716 22596 30772 22606
rect 30492 22372 30548 22382
rect 30492 22278 30548 22316
rect 30268 22194 30324 22204
rect 30604 22260 30660 22270
rect 30716 22260 30772 22540
rect 30660 22204 30772 22260
rect 30604 22194 30660 22204
rect 30156 21476 30212 21486
rect 29932 20862 29934 20914
rect 29986 20862 29988 20914
rect 29484 20580 29540 20590
rect 29484 20486 29540 20524
rect 29148 20132 29316 20188
rect 28700 19906 28756 19918
rect 28700 19854 28702 19906
rect 28754 19854 28756 19906
rect 28700 19794 28756 19854
rect 28700 19742 28702 19794
rect 28754 19742 28756 19794
rect 28700 19730 28756 19742
rect 28588 19684 28644 19694
rect 28588 19346 28644 19628
rect 29148 19684 29204 20132
rect 29260 19908 29316 19918
rect 29260 19906 29428 19908
rect 29260 19854 29262 19906
rect 29314 19854 29428 19906
rect 29260 19852 29428 19854
rect 29260 19842 29316 19852
rect 29148 19618 29204 19628
rect 28588 19294 28590 19346
rect 28642 19294 28644 19346
rect 28588 18564 28644 19294
rect 28588 18498 28644 18508
rect 29148 19348 29204 19358
rect 28924 18338 28980 18350
rect 28924 18286 28926 18338
rect 28978 18286 28980 18338
rect 28476 16930 28532 16940
rect 28588 18116 28644 18126
rect 28588 17778 28644 18060
rect 28924 18116 28980 18286
rect 28924 18050 28980 18060
rect 28588 17726 28590 17778
rect 28642 17726 28644 17778
rect 28364 16818 28420 16828
rect 28476 16772 28532 16782
rect 28252 16370 28308 16380
rect 28364 16548 28420 16558
rect 28364 16210 28420 16492
rect 28364 16158 28366 16210
rect 28418 16158 28420 16210
rect 28364 16146 28420 16158
rect 28140 15314 28196 15484
rect 28140 15262 28142 15314
rect 28194 15262 28196 15314
rect 28140 15250 28196 15262
rect 28252 16100 28308 16110
rect 28252 15148 28308 16044
rect 28028 15026 28084 15036
rect 28140 15092 28308 15148
rect 28364 15988 28420 15998
rect 27916 14644 27972 14654
rect 28140 14644 28196 15092
rect 27916 14642 28196 14644
rect 27916 14590 27918 14642
rect 27970 14590 28196 14642
rect 27916 14588 28196 14590
rect 27916 14578 27972 14588
rect 28028 14308 28084 14318
rect 28028 13746 28084 14252
rect 28028 13694 28030 13746
rect 28082 13694 28084 13746
rect 28028 13636 28084 13694
rect 28028 13570 28084 13580
rect 27468 13468 27636 13524
rect 26908 12178 27300 12180
rect 26908 12126 26910 12178
rect 26962 12126 27300 12178
rect 26908 12124 27300 12126
rect 27356 13076 27412 13086
rect 27356 12178 27412 13020
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 26908 12114 26964 12124
rect 27356 12114 27412 12126
rect 26460 11954 26516 11966
rect 27132 11956 27188 11966
rect 26460 11902 26462 11954
rect 26514 11902 26516 11954
rect 26348 10164 26404 10174
rect 26348 9604 26404 10108
rect 26460 9828 26516 11902
rect 27020 11900 27132 11956
rect 26908 11732 26964 11742
rect 26684 11620 26740 11630
rect 26684 10834 26740 11564
rect 26908 11394 26964 11676
rect 26908 11342 26910 11394
rect 26962 11342 26964 11394
rect 26908 11330 26964 11342
rect 26684 10782 26686 10834
rect 26738 10782 26740 10834
rect 26572 10724 26628 10734
rect 26572 10630 26628 10668
rect 26684 10052 26740 10782
rect 26684 9986 26740 9996
rect 26796 10276 26852 10286
rect 26684 9828 26740 9838
rect 26460 9826 26740 9828
rect 26460 9774 26686 9826
rect 26738 9774 26740 9826
rect 26460 9772 26740 9774
rect 26684 9762 26740 9772
rect 26460 9604 26516 9614
rect 26348 9602 26516 9604
rect 26348 9550 26462 9602
rect 26514 9550 26516 9602
rect 26348 9548 26516 9550
rect 26460 9538 26516 9548
rect 26572 9604 26628 9614
rect 26796 9604 26852 10220
rect 26572 9602 26852 9604
rect 26572 9550 26574 9602
rect 26626 9550 26852 9602
rect 26572 9548 26852 9550
rect 26572 9538 26628 9548
rect 26684 9380 26740 9390
rect 26684 9154 26740 9324
rect 26908 9268 26964 9278
rect 27020 9268 27076 11900
rect 27132 11862 27188 11900
rect 27468 11732 27524 13468
rect 28364 13412 28420 15932
rect 28476 15874 28532 16716
rect 28588 16100 28644 17726
rect 28924 16772 28980 16782
rect 28588 16034 28644 16044
rect 28700 16100 28756 16110
rect 28924 16100 28980 16716
rect 28700 16098 28980 16100
rect 28700 16046 28702 16098
rect 28754 16046 28980 16098
rect 28700 16044 28980 16046
rect 28700 16034 28756 16044
rect 28476 15822 28478 15874
rect 28530 15822 28532 15874
rect 28476 15764 28532 15822
rect 28476 15698 28532 15708
rect 28588 15428 28644 15438
rect 28476 15314 28532 15326
rect 28476 15262 28478 15314
rect 28530 15262 28532 15314
rect 28476 15092 28532 15262
rect 28476 15026 28532 15036
rect 28476 14868 28532 14878
rect 28476 13860 28532 14812
rect 28588 14532 28644 15372
rect 28700 15426 28756 15438
rect 28700 15374 28702 15426
rect 28754 15374 28756 15426
rect 28700 14756 28756 15374
rect 28812 15204 28868 15214
rect 28812 15110 28868 15148
rect 28700 14690 28756 14700
rect 28588 14466 28644 14476
rect 28812 14420 28868 14430
rect 28812 14326 28868 14364
rect 28588 14306 28644 14318
rect 28588 14254 28590 14306
rect 28642 14254 28644 14306
rect 28588 14084 28644 14254
rect 28588 14018 28644 14028
rect 28700 14306 28756 14318
rect 28700 14254 28702 14306
rect 28754 14254 28756 14306
rect 28476 13728 28532 13804
rect 28364 13346 28420 13356
rect 28588 13412 28644 13422
rect 28252 13300 28308 13310
rect 27804 13186 27860 13198
rect 27804 13134 27806 13186
rect 27858 13134 27860 13186
rect 27692 12852 27748 12862
rect 27692 12758 27748 12796
rect 27468 11666 27524 11676
rect 27580 12292 27636 12302
rect 27244 11284 27300 11294
rect 27244 9492 27300 11228
rect 27580 11060 27636 12236
rect 27580 10994 27636 11004
rect 27468 10612 27524 10622
rect 27468 10610 27636 10612
rect 27468 10558 27470 10610
rect 27522 10558 27636 10610
rect 27468 10556 27636 10558
rect 27468 10546 27524 10556
rect 27356 9828 27412 9838
rect 27356 9734 27412 9772
rect 27468 9716 27524 9726
rect 27468 9622 27524 9660
rect 27580 9492 27636 10556
rect 27804 10164 27860 13134
rect 27916 12740 27972 12750
rect 28140 12740 28196 12750
rect 27916 12738 28084 12740
rect 27916 12686 27918 12738
rect 27970 12686 28084 12738
rect 27916 12684 28084 12686
rect 27916 12674 27972 12684
rect 27916 11956 27972 11966
rect 27916 11284 27972 11900
rect 27916 11218 27972 11228
rect 27916 10836 27972 10846
rect 28028 10836 28084 12684
rect 28140 12646 28196 12684
rect 28252 12292 28308 13244
rect 28476 13188 28532 13198
rect 28364 12852 28420 12862
rect 28364 12758 28420 12796
rect 28252 12198 28308 12236
rect 28364 12178 28420 12190
rect 28364 12126 28366 12178
rect 28418 12126 28420 12178
rect 28252 11956 28308 11966
rect 28252 11862 28308 11900
rect 28364 10948 28420 12126
rect 28476 11956 28532 13132
rect 28476 11890 28532 11900
rect 28588 12740 28644 13356
rect 28700 12964 28756 14254
rect 28700 12898 28756 12908
rect 28924 14308 28980 16044
rect 29148 14756 29204 19292
rect 29372 19012 29428 19852
rect 29596 19906 29652 19918
rect 29596 19854 29598 19906
rect 29650 19854 29652 19906
rect 29036 14700 29204 14756
rect 29260 18228 29316 18238
rect 29036 14644 29092 14700
rect 29036 14578 29092 14588
rect 28812 12740 28868 12750
rect 28588 12738 28868 12740
rect 28588 12686 28814 12738
rect 28866 12686 28868 12738
rect 28588 12684 28868 12686
rect 28588 11732 28644 12684
rect 28812 12674 28868 12684
rect 28924 12290 28980 14252
rect 29148 14532 29204 14542
rect 29260 14532 29316 18172
rect 29372 18116 29428 18956
rect 29484 19794 29540 19806
rect 29484 19742 29486 19794
rect 29538 19742 29540 19794
rect 29484 19010 29540 19742
rect 29596 19236 29652 19854
rect 29932 19348 29988 20862
rect 30044 21474 30212 21476
rect 30044 21422 30158 21474
rect 30210 21422 30212 21474
rect 30044 21420 30212 21422
rect 30044 19796 30100 21420
rect 30156 21410 30212 21420
rect 30492 21476 30548 21486
rect 30492 21474 30660 21476
rect 30492 21422 30494 21474
rect 30546 21422 30660 21474
rect 30492 21420 30660 21422
rect 30492 21410 30548 21420
rect 30492 20578 30548 20590
rect 30492 20526 30494 20578
rect 30546 20526 30548 20578
rect 30156 19908 30212 19918
rect 30156 19814 30212 19852
rect 30492 19906 30548 20526
rect 30604 20244 30660 21420
rect 30716 20356 30772 22204
rect 30716 20290 30772 20300
rect 30604 20178 30660 20188
rect 30492 19854 30494 19906
rect 30546 19854 30548 19906
rect 30044 19730 30100 19740
rect 29932 19282 29988 19292
rect 29596 19170 29652 19180
rect 29484 18958 29486 19010
rect 29538 18958 29540 19010
rect 29484 18452 29540 18958
rect 29932 19012 29988 19022
rect 30492 19012 30548 19854
rect 30828 19796 30884 22990
rect 31388 22708 31444 22718
rect 31388 22482 31444 22652
rect 31500 22596 31556 23662
rect 31724 23268 31780 23278
rect 31500 22530 31556 22540
rect 31612 23042 31668 23054
rect 31612 22990 31614 23042
rect 31666 22990 31668 23042
rect 31388 22430 31390 22482
rect 31442 22430 31444 22482
rect 31388 22418 31444 22430
rect 30940 22146 30996 22158
rect 30940 22094 30942 22146
rect 30994 22094 30996 22146
rect 30940 21924 30996 22094
rect 30940 21858 30996 21868
rect 31276 22148 31332 22158
rect 31276 21700 31332 22092
rect 31612 21812 31668 22990
rect 31612 21746 31668 21756
rect 31724 22482 31780 23212
rect 31836 23156 31892 24558
rect 31836 23090 31892 23100
rect 32060 24162 32116 24174
rect 32060 24110 32062 24162
rect 32114 24110 32116 24162
rect 32060 23714 32116 24110
rect 32956 24162 33012 24174
rect 32956 24110 32958 24162
rect 33010 24110 33012 24162
rect 32956 24050 33012 24110
rect 32956 23998 32958 24050
rect 33010 23998 33012 24050
rect 32956 23986 33012 23998
rect 33068 23828 33124 25228
rect 35756 24724 35812 24734
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35756 24052 35812 24668
rect 34188 23940 34244 23950
rect 35756 23920 35812 23996
rect 35980 24612 36036 24622
rect 34188 23846 34244 23884
rect 32956 23772 33124 23828
rect 32060 23662 32062 23714
rect 32114 23662 32116 23714
rect 31724 22430 31726 22482
rect 31778 22430 31780 22482
rect 31052 21474 31108 21486
rect 31052 21422 31054 21474
rect 31106 21422 31108 21474
rect 30828 19730 30884 19740
rect 30940 20578 30996 20590
rect 30940 20526 30942 20578
rect 30994 20526 30996 20578
rect 30716 19012 30772 19022
rect 30492 19010 30772 19012
rect 30492 18958 30718 19010
rect 30770 18958 30772 19010
rect 30492 18956 30772 18958
rect 29932 18918 29988 18956
rect 30716 18900 30772 18956
rect 29820 18676 29876 18686
rect 29484 18386 29540 18396
rect 29596 18674 29876 18676
rect 29596 18622 29822 18674
rect 29874 18622 29876 18674
rect 29596 18620 29876 18622
rect 29372 18050 29428 18060
rect 29596 16548 29652 18620
rect 29820 18610 29876 18620
rect 29596 16482 29652 16492
rect 29708 18452 29764 18462
rect 29484 15874 29540 15886
rect 29484 15822 29486 15874
rect 29538 15822 29540 15874
rect 29484 15652 29540 15822
rect 29484 15586 29540 15596
rect 29596 15874 29652 15886
rect 29596 15822 29598 15874
rect 29650 15822 29652 15874
rect 29596 15540 29652 15822
rect 29708 15540 29764 18396
rect 29932 18450 29988 18462
rect 29932 18398 29934 18450
rect 29986 18398 29988 18450
rect 29932 18340 29988 18398
rect 30604 18340 30660 18350
rect 30716 18340 30772 18844
rect 30940 18564 30996 20526
rect 31052 20188 31108 21422
rect 31276 20914 31332 21644
rect 31724 21700 31780 22430
rect 31948 23042 32004 23054
rect 31948 22990 31950 23042
rect 32002 22990 32004 23042
rect 31724 21634 31780 21644
rect 31836 22260 31892 22270
rect 31724 21476 31780 21486
rect 31836 21476 31892 22204
rect 31780 21420 31892 21476
rect 31724 21382 31780 21420
rect 31276 20862 31278 20914
rect 31330 20862 31332 20914
rect 31276 20850 31332 20862
rect 31836 20580 31892 20590
rect 31836 20486 31892 20524
rect 31836 20244 31892 20254
rect 31052 20132 31332 20188
rect 31836 20150 31892 20188
rect 31052 19908 31108 19918
rect 31052 19012 31108 19852
rect 31052 18946 31108 18956
rect 31164 19010 31220 19022
rect 31164 18958 31166 19010
rect 31218 18958 31220 19010
rect 30940 18498 30996 18508
rect 29932 18284 30436 18340
rect 29820 18228 29876 18238
rect 29820 18226 29988 18228
rect 29820 18174 29822 18226
rect 29874 18174 29988 18226
rect 29820 18172 29988 18174
rect 29820 18162 29876 18172
rect 29820 17442 29876 17454
rect 29820 17390 29822 17442
rect 29874 17390 29876 17442
rect 29820 17220 29876 17390
rect 29820 17154 29876 17164
rect 29932 16996 29988 18172
rect 30044 18116 30100 18126
rect 30044 17666 30100 18060
rect 30044 17614 30046 17666
rect 30098 17614 30100 17666
rect 30044 17602 30100 17614
rect 30268 17668 30324 17678
rect 30268 17574 30324 17612
rect 30156 17444 30212 17454
rect 30156 17350 30212 17388
rect 29820 16940 29988 16996
rect 30380 16996 30436 18284
rect 30660 18284 30772 18340
rect 31052 18340 31108 18350
rect 30492 18228 30548 18238
rect 30492 18134 30548 18172
rect 29820 16548 29876 16940
rect 30380 16884 30436 16940
rect 30156 16882 30436 16884
rect 30156 16830 30382 16882
rect 30434 16830 30436 16882
rect 30156 16828 30436 16830
rect 29932 16772 29988 16782
rect 29932 16678 29988 16716
rect 30044 16548 30100 16558
rect 29820 16492 29988 16548
rect 29820 15876 29876 15886
rect 29820 15782 29876 15820
rect 29708 15484 29876 15540
rect 29596 15474 29652 15484
rect 29484 15428 29540 15438
rect 29372 15316 29428 15326
rect 29372 15222 29428 15260
rect 29484 15204 29540 15372
rect 29708 15316 29764 15326
rect 29708 15222 29764 15260
rect 29484 15138 29540 15148
rect 29596 14532 29652 14542
rect 29260 14530 29652 14532
rect 29260 14478 29598 14530
rect 29650 14478 29652 14530
rect 29260 14476 29652 14478
rect 28924 12238 28926 12290
rect 28978 12238 28980 12290
rect 28924 12226 28980 12238
rect 29036 14196 29092 14206
rect 28364 10882 28420 10892
rect 28476 11676 28644 11732
rect 28028 10780 28196 10836
rect 27916 10722 27972 10780
rect 27916 10670 27918 10722
rect 27970 10670 27972 10722
rect 27916 10658 27972 10670
rect 27804 10098 27860 10108
rect 28028 10612 28084 10622
rect 27692 9940 27748 9950
rect 27692 9846 27748 9884
rect 27244 9436 27412 9492
rect 26908 9266 27076 9268
rect 26908 9214 26910 9266
rect 26962 9214 27076 9266
rect 26908 9212 27076 9214
rect 27132 9380 27188 9390
rect 27132 9266 27188 9324
rect 27132 9214 27134 9266
rect 27186 9214 27188 9266
rect 26908 9202 26964 9212
rect 27132 9202 27188 9214
rect 27244 9268 27300 9278
rect 27244 9174 27300 9212
rect 26684 9102 26686 9154
rect 26738 9102 26740 9154
rect 26684 9090 26740 9102
rect 26236 7586 26292 8764
rect 26796 8596 26852 8606
rect 26236 7534 26238 7586
rect 26290 7534 26292 7586
rect 26236 7522 26292 7534
rect 26460 8036 26516 8046
rect 25676 6638 25678 6690
rect 25730 6638 25732 6690
rect 25676 6626 25732 6638
rect 25788 7476 25844 7486
rect 25004 5294 25006 5346
rect 25058 5294 25060 5346
rect 25004 5282 25060 5294
rect 25228 6580 25284 6590
rect 25228 5124 25284 6524
rect 25564 6468 25620 6478
rect 25788 6468 25844 7420
rect 26460 7474 26516 7980
rect 26796 7698 26852 8540
rect 26796 7646 26798 7698
rect 26850 7646 26852 7698
rect 26796 7634 26852 7646
rect 26908 7812 26964 7822
rect 26460 7422 26462 7474
rect 26514 7422 26516 7474
rect 26460 7410 26516 7422
rect 25564 6374 25620 6412
rect 25676 6412 25844 6468
rect 25900 6690 25956 6702
rect 25900 6638 25902 6690
rect 25954 6638 25956 6690
rect 25564 6132 25620 6142
rect 25564 6038 25620 6076
rect 25228 5058 25284 5068
rect 25340 5684 25396 5694
rect 24780 5012 24836 5022
rect 24780 4562 24836 4956
rect 24780 4510 24782 4562
rect 24834 4510 24836 4562
rect 24780 4498 24836 4510
rect 24892 5010 24948 5022
rect 24892 4958 24894 5010
rect 24946 4958 24948 5010
rect 24892 4564 24948 4958
rect 24948 4508 25060 4564
rect 24892 4498 24948 4508
rect 24892 4338 24948 4350
rect 24892 4286 24894 4338
rect 24946 4286 24948 4338
rect 24892 4228 24948 4286
rect 24556 3332 24724 3388
rect 24668 2884 24724 3332
rect 24668 2818 24724 2828
rect 24892 2772 24948 4172
rect 25004 3444 25060 4508
rect 25340 3666 25396 5628
rect 25564 5236 25620 5246
rect 25564 5142 25620 5180
rect 25340 3614 25342 3666
rect 25394 3614 25396 3666
rect 25340 3602 25396 3614
rect 25452 4452 25508 4462
rect 25004 3332 25060 3388
rect 25004 3266 25060 3276
rect 25452 3220 25508 4396
rect 25676 4450 25732 6412
rect 25900 6132 25956 6638
rect 26348 6690 26404 6702
rect 26348 6638 26350 6690
rect 26402 6638 26404 6690
rect 26348 6356 26404 6638
rect 26796 6578 26852 6590
rect 26796 6526 26798 6578
rect 26850 6526 26852 6578
rect 26348 6290 26404 6300
rect 26684 6466 26740 6478
rect 26684 6414 26686 6466
rect 26738 6414 26740 6466
rect 26012 6132 26068 6142
rect 25900 6130 26068 6132
rect 25900 6078 26014 6130
rect 26066 6078 26068 6130
rect 25900 6076 26068 6078
rect 26012 6066 26068 6076
rect 25788 5908 25844 5918
rect 25788 4562 25844 5852
rect 26124 5906 26180 5918
rect 26124 5854 26126 5906
rect 26178 5854 26180 5906
rect 26124 5796 26180 5854
rect 26348 5908 26404 5918
rect 26348 5814 26404 5852
rect 26684 5908 26740 6414
rect 26796 6132 26852 6526
rect 26908 6468 26964 7756
rect 27020 6692 27076 6702
rect 27020 6598 27076 6636
rect 27132 6580 27188 6590
rect 26908 6412 27076 6468
rect 26796 6076 26964 6132
rect 26684 5842 26740 5852
rect 26796 5906 26852 5918
rect 26796 5854 26798 5906
rect 26850 5854 26852 5906
rect 26124 5348 26180 5740
rect 26572 5682 26628 5694
rect 26572 5630 26574 5682
rect 26626 5630 26628 5682
rect 26572 5572 26628 5630
rect 26572 5506 26628 5516
rect 26796 5460 26852 5854
rect 26796 5394 26852 5404
rect 26124 5282 26180 5292
rect 26572 5010 26628 5022
rect 26572 4958 26574 5010
rect 26626 4958 26628 5010
rect 25788 4510 25790 4562
rect 25842 4510 25844 4562
rect 25788 4498 25844 4510
rect 26012 4564 26068 4574
rect 26012 4470 26068 4508
rect 25676 4398 25678 4450
rect 25730 4398 25732 4450
rect 25676 4386 25732 4398
rect 26572 4452 26628 4958
rect 26572 4386 26628 4396
rect 26908 5012 26964 6076
rect 27020 6018 27076 6412
rect 27020 5966 27022 6018
rect 27074 5966 27076 6018
rect 27020 5572 27076 5966
rect 27020 5506 27076 5516
rect 26460 4340 26516 4350
rect 26460 4246 26516 4284
rect 26348 3780 26404 3790
rect 24892 2706 24948 2716
rect 25340 3164 25508 3220
rect 25788 3444 25844 3454
rect 25340 800 25396 3164
rect 25788 1652 25844 3388
rect 26348 3442 26404 3724
rect 26908 3556 26964 4956
rect 27132 5236 27188 6524
rect 27356 6020 27412 9436
rect 27468 9436 27636 9492
rect 27804 9714 27860 9726
rect 27804 9662 27806 9714
rect 27858 9662 27860 9714
rect 27468 7812 27524 9436
rect 27804 9380 27860 9662
rect 27468 7746 27524 7756
rect 27580 9324 27860 9380
rect 27356 5954 27412 5964
rect 27468 7474 27524 7486
rect 27468 7422 27470 7474
rect 27522 7422 27524 7474
rect 27132 3556 27188 5180
rect 27468 5460 27524 7422
rect 27580 6132 27636 9324
rect 27804 9156 27860 9166
rect 27804 9062 27860 9100
rect 27916 9044 27972 9054
rect 27916 8950 27972 8988
rect 27804 8820 27860 8830
rect 28028 8820 28084 10556
rect 28140 9828 28196 10780
rect 28364 10724 28420 10734
rect 28364 10630 28420 10668
rect 28140 9762 28196 9772
rect 28252 9602 28308 9614
rect 28252 9550 28254 9602
rect 28306 9550 28308 9602
rect 28252 8932 28308 9550
rect 28252 8866 28308 8876
rect 28364 9602 28420 9614
rect 28364 9550 28366 9602
rect 28418 9550 28420 9602
rect 27804 8818 28084 8820
rect 27804 8766 27806 8818
rect 27858 8766 28084 8818
rect 27804 8764 28084 8766
rect 27804 8754 27860 8764
rect 28364 8596 28420 9550
rect 28476 9268 28532 11676
rect 28700 11508 28756 11518
rect 28924 11508 28980 11518
rect 28700 11414 28756 11452
rect 28812 11452 28924 11508
rect 28700 11060 28756 11070
rect 28588 10722 28644 10734
rect 28588 10670 28590 10722
rect 28642 10670 28644 10722
rect 28588 9828 28644 10670
rect 28700 10610 28756 11004
rect 28700 10558 28702 10610
rect 28754 10558 28756 10610
rect 28700 10388 28756 10558
rect 28700 10322 28756 10332
rect 28588 9772 28756 9828
rect 28588 9604 28644 9614
rect 28588 9510 28644 9548
rect 28476 9202 28532 9212
rect 28588 9156 28644 9166
rect 28588 9062 28644 9100
rect 28364 8530 28420 8540
rect 28476 9042 28532 9054
rect 28476 8990 28478 9042
rect 28530 8990 28532 9042
rect 28476 7700 28532 8990
rect 28700 8370 28756 9772
rect 28812 9826 28868 11452
rect 28924 11442 28980 11452
rect 28812 9774 28814 9826
rect 28866 9774 28868 9826
rect 28812 9716 28868 9774
rect 28812 9650 28868 9660
rect 28924 10052 28980 10062
rect 28700 8318 28702 8370
rect 28754 8318 28756 8370
rect 28700 7924 28756 8318
rect 28700 7858 28756 7868
rect 28812 9042 28868 9054
rect 28812 8990 28814 9042
rect 28866 8990 28868 9042
rect 28812 7700 28868 8990
rect 28364 7644 28532 7700
rect 28700 7644 28868 7700
rect 27916 7588 27972 7598
rect 27692 7364 27748 7374
rect 27692 6578 27748 7308
rect 27916 7140 27972 7532
rect 27916 7074 27972 7084
rect 28140 7476 28196 7486
rect 28140 6690 28196 7420
rect 28140 6638 28142 6690
rect 28194 6638 28196 6690
rect 28140 6626 28196 6638
rect 27692 6526 27694 6578
rect 27746 6526 27748 6578
rect 27692 6514 27748 6526
rect 27916 6468 27972 6478
rect 27916 6374 27972 6412
rect 28028 6466 28084 6478
rect 28028 6414 28030 6466
rect 28082 6414 28084 6466
rect 27692 6132 27748 6142
rect 27580 6130 27748 6132
rect 27580 6078 27694 6130
rect 27746 6078 27748 6130
rect 27580 6076 27748 6078
rect 27692 6066 27748 6076
rect 27580 5908 27636 5918
rect 27580 5814 27636 5852
rect 27468 5124 27524 5404
rect 27468 5058 27524 5068
rect 27804 5572 27860 5582
rect 27804 5122 27860 5516
rect 27804 5070 27806 5122
rect 27858 5070 27860 5122
rect 27804 5058 27860 5070
rect 28028 4788 28084 6414
rect 28364 5908 28420 7644
rect 28476 7476 28532 7486
rect 28476 7382 28532 7420
rect 28588 7364 28644 7374
rect 28588 7270 28644 7308
rect 28700 6690 28756 7644
rect 28812 7474 28868 7486
rect 28812 7422 28814 7474
rect 28866 7422 28868 7474
rect 28812 7364 28868 7422
rect 28812 7298 28868 7308
rect 28700 6638 28702 6690
rect 28754 6638 28756 6690
rect 28700 6626 28756 6638
rect 28812 7140 28868 7150
rect 28812 6690 28868 7084
rect 28812 6638 28814 6690
rect 28866 6638 28868 6690
rect 28812 6626 28868 6638
rect 28364 5842 28420 5852
rect 28476 6020 28532 6030
rect 28252 5796 28308 5806
rect 28252 5702 28308 5740
rect 28364 5348 28420 5358
rect 28364 5254 28420 5292
rect 27804 4732 28084 4788
rect 28140 5010 28196 5022
rect 28140 4958 28142 5010
rect 28194 4958 28196 5010
rect 27244 4228 27300 4238
rect 27244 4226 27748 4228
rect 27244 4174 27246 4226
rect 27298 4174 27748 4226
rect 27244 4172 27748 4174
rect 27244 4162 27300 4172
rect 27692 3666 27748 4172
rect 27692 3614 27694 3666
rect 27746 3614 27748 3666
rect 27692 3602 27748 3614
rect 27356 3556 27412 3566
rect 27132 3554 27412 3556
rect 27132 3502 27358 3554
rect 27410 3502 27412 3554
rect 27132 3500 27412 3502
rect 26908 3490 26964 3500
rect 27356 3490 27412 3500
rect 27580 3556 27636 3566
rect 27580 3462 27636 3500
rect 27804 3554 27860 4732
rect 28140 4564 28196 4958
rect 28140 4498 28196 4508
rect 28252 4898 28308 4910
rect 28252 4846 28254 4898
rect 28306 4846 28308 4898
rect 28252 4228 28308 4846
rect 27804 3502 27806 3554
rect 27858 3502 27860 3554
rect 27804 3490 27860 3502
rect 28028 4172 28308 4228
rect 28028 3554 28084 4172
rect 28028 3502 28030 3554
rect 28082 3502 28084 3554
rect 28028 3490 28084 3502
rect 26348 3390 26350 3442
rect 26402 3390 26404 3442
rect 26348 3378 26404 3390
rect 26684 3444 26740 3454
rect 28476 3388 28532 5964
rect 28588 5460 28644 5470
rect 28588 5234 28644 5404
rect 28588 5182 28590 5234
rect 28642 5182 28644 5234
rect 28588 5170 28644 5182
rect 28812 5236 28868 5246
rect 28812 5122 28868 5180
rect 28812 5070 28814 5122
rect 28866 5070 28868 5122
rect 28812 5058 28868 5070
rect 28588 3668 28644 3678
rect 28924 3668 28980 9996
rect 29036 9154 29092 14140
rect 29148 13188 29204 14476
rect 29596 14466 29652 14476
rect 29708 14532 29764 14542
rect 29708 14418 29764 14476
rect 29708 14366 29710 14418
rect 29762 14366 29764 14418
rect 29708 14354 29764 14366
rect 29596 14084 29652 14094
rect 29260 13746 29316 13758
rect 29260 13694 29262 13746
rect 29314 13694 29316 13746
rect 29260 13524 29316 13694
rect 29260 13458 29316 13468
rect 29372 13636 29428 13646
rect 29148 13132 29316 13188
rect 29148 12180 29204 12190
rect 29148 10836 29204 12124
rect 29148 10770 29204 10780
rect 29260 11956 29316 13132
rect 29372 12180 29428 13580
rect 29484 12962 29540 12974
rect 29484 12910 29486 12962
rect 29538 12910 29540 12962
rect 29484 12402 29540 12910
rect 29596 12852 29652 14028
rect 29820 13524 29876 15484
rect 29932 15426 29988 16492
rect 29932 15374 29934 15426
rect 29986 15374 29988 15426
rect 29932 15362 29988 15374
rect 30044 15876 30100 16492
rect 30156 16098 30212 16828
rect 30380 16818 30436 16828
rect 30492 18004 30548 18014
rect 30492 16436 30548 17948
rect 30604 17220 30660 18284
rect 31052 18246 31108 18284
rect 31164 18116 31220 18958
rect 31164 18050 31220 18060
rect 30940 17780 30996 17790
rect 30940 17686 30996 17724
rect 31276 17780 31332 20132
rect 31388 19906 31444 19918
rect 31388 19854 31390 19906
rect 31442 19854 31444 19906
rect 31388 19796 31444 19854
rect 31388 19730 31444 19740
rect 31948 19684 32004 22990
rect 32060 19908 32116 23662
rect 32508 23714 32564 23726
rect 32508 23662 32510 23714
rect 32562 23662 32564 23714
rect 32508 23604 32564 23662
rect 32508 23538 32564 23548
rect 32956 23378 33012 23772
rect 33292 23716 33348 23726
rect 33292 23622 33348 23660
rect 33852 23714 33908 23726
rect 33852 23662 33854 23714
rect 33906 23662 33908 23714
rect 32956 23326 32958 23378
rect 33010 23326 33012 23378
rect 32956 23314 33012 23326
rect 32172 23268 32228 23278
rect 32172 22482 32228 23212
rect 32508 23268 32564 23278
rect 32508 23174 32564 23212
rect 33404 23268 33460 23278
rect 32172 22430 32174 22482
rect 32226 22430 32228 22482
rect 32172 22418 32228 22430
rect 32620 23044 32676 23054
rect 32620 22482 32676 22988
rect 32620 22430 32622 22482
rect 32674 22430 32676 22482
rect 32620 22418 32676 22430
rect 32508 22372 32564 22382
rect 33404 22372 33460 23212
rect 33516 23044 33572 23054
rect 33516 22950 33572 22988
rect 33852 23044 33908 23662
rect 35308 23716 35364 23726
rect 35308 23622 35364 23660
rect 35084 23156 35140 23166
rect 33852 22978 33908 22988
rect 33964 23042 34020 23054
rect 33964 22990 33966 23042
rect 34018 22990 34020 23042
rect 33964 22932 34020 22990
rect 33964 22866 34020 22876
rect 34188 23044 34244 23054
rect 34188 22482 34244 22988
rect 34188 22430 34190 22482
rect 34242 22430 34244 22482
rect 34188 22418 34244 22430
rect 34524 23042 34580 23054
rect 34524 22990 34526 23042
rect 34578 22990 34580 23042
rect 33404 22316 33572 22372
rect 32172 21812 32228 21822
rect 32172 21718 32228 21756
rect 32284 20578 32340 20590
rect 32284 20526 32286 20578
rect 32338 20526 32340 20578
rect 32284 20188 32340 20526
rect 32284 20132 32452 20188
rect 32060 19842 32116 19852
rect 32284 19906 32340 19918
rect 32284 19854 32286 19906
rect 32338 19854 32340 19906
rect 31276 17714 31332 17724
rect 31500 19012 31556 19022
rect 31500 18338 31556 18956
rect 31612 19010 31668 19022
rect 31612 18958 31614 19010
rect 31666 18958 31668 19010
rect 31612 18900 31668 18958
rect 31612 18834 31668 18844
rect 31948 18788 32004 19628
rect 32284 19460 32340 19854
rect 32284 19394 32340 19404
rect 31948 18722 32004 18732
rect 32284 19236 32340 19246
rect 32284 19010 32340 19180
rect 32284 18958 32286 19010
rect 32338 18958 32340 19010
rect 31500 18286 31502 18338
rect 31554 18286 31556 18338
rect 31500 17668 31556 18286
rect 31948 18338 32004 18350
rect 31948 18286 31950 18338
rect 32002 18286 32004 18338
rect 31948 18116 32004 18286
rect 31948 18050 32004 18060
rect 31500 17602 31556 17612
rect 31612 18004 31668 18014
rect 31052 17556 31108 17566
rect 31052 17462 31108 17500
rect 30604 17154 30660 17164
rect 30828 17442 30884 17454
rect 30828 17390 30830 17442
rect 30882 17390 30884 17442
rect 30716 16882 30772 16894
rect 30716 16830 30718 16882
rect 30770 16830 30772 16882
rect 30716 16548 30772 16830
rect 30828 16770 30884 17390
rect 31276 17444 31332 17454
rect 31276 17350 31332 17388
rect 31500 17444 31556 17454
rect 30828 16718 30830 16770
rect 30882 16718 30884 16770
rect 30828 16706 30884 16718
rect 30940 16994 30996 17006
rect 30940 16942 30942 16994
rect 30994 16942 30996 16994
rect 30716 16482 30772 16492
rect 30492 16380 30660 16436
rect 30604 16212 30660 16380
rect 30716 16212 30772 16222
rect 30604 16210 30772 16212
rect 30604 16158 30718 16210
rect 30770 16158 30772 16210
rect 30604 16156 30772 16158
rect 30716 16146 30772 16156
rect 30156 16046 30158 16098
rect 30210 16046 30212 16098
rect 30156 16034 30212 16046
rect 30940 16100 30996 16942
rect 31388 16996 31444 17006
rect 31388 16902 31444 16940
rect 30940 16034 30996 16044
rect 31276 16660 31332 16670
rect 31276 16098 31332 16604
rect 31500 16212 31556 17388
rect 31612 17106 31668 17948
rect 31836 17444 31892 17454
rect 31612 17054 31614 17106
rect 31666 17054 31668 17106
rect 31612 17042 31668 17054
rect 31724 17442 31892 17444
rect 31724 17390 31838 17442
rect 31890 17390 31892 17442
rect 31724 17388 31892 17390
rect 31724 17220 31780 17388
rect 31836 17378 31892 17388
rect 31724 16994 31780 17164
rect 31724 16942 31726 16994
rect 31778 16942 31780 16994
rect 31724 16930 31780 16942
rect 32060 17220 32116 17230
rect 31724 16660 31780 16670
rect 31500 16156 31668 16212
rect 31276 16046 31278 16098
rect 31330 16046 31332 16098
rect 31276 16034 31332 16046
rect 31500 15988 31556 15998
rect 30604 15876 30660 15886
rect 30044 15148 30100 15820
rect 30492 15874 30660 15876
rect 30492 15822 30606 15874
rect 30658 15822 30660 15874
rect 30492 15820 30660 15822
rect 29932 15092 30100 15148
rect 30156 15764 30212 15774
rect 29932 14306 29988 15092
rect 29932 14254 29934 14306
rect 29986 14254 29988 14306
rect 29932 13860 29988 14254
rect 29932 13794 29988 13804
rect 29820 13458 29876 13468
rect 29932 13634 29988 13646
rect 29932 13582 29934 13634
rect 29986 13582 29988 13634
rect 29708 13076 29764 13086
rect 29932 13076 29988 13582
rect 30156 13188 30212 15708
rect 30380 15540 30436 15550
rect 30380 15446 30436 15484
rect 30268 15316 30324 15326
rect 30268 14530 30324 15260
rect 30268 14478 30270 14530
rect 30322 14478 30324 14530
rect 30268 14466 30324 14478
rect 30492 14532 30548 15820
rect 30604 15810 30660 15820
rect 31388 15874 31444 15886
rect 31388 15822 31390 15874
rect 31442 15822 31444 15874
rect 30604 15540 30660 15550
rect 30604 15446 30660 15484
rect 31388 15540 31444 15822
rect 31388 15474 31444 15484
rect 31500 15538 31556 15932
rect 31500 15486 31502 15538
rect 31554 15486 31556 15538
rect 31500 15474 31556 15486
rect 31612 15538 31668 16156
rect 31612 15486 31614 15538
rect 31666 15486 31668 15538
rect 30716 15316 30772 15326
rect 30716 15222 30772 15260
rect 31500 15204 31556 15214
rect 31388 15092 31556 15148
rect 30492 14466 30548 14476
rect 30828 14868 30884 14878
rect 30604 14420 30660 14430
rect 30604 14326 30660 14364
rect 30492 14308 30548 14318
rect 30492 14214 30548 14252
rect 29708 13074 29988 13076
rect 29708 13022 29710 13074
rect 29762 13022 29988 13074
rect 29708 13020 29988 13022
rect 30044 13132 30212 13188
rect 30492 13860 30548 13870
rect 29708 13010 29764 13020
rect 29932 12852 29988 12862
rect 30044 12852 30100 13132
rect 30156 12964 30212 12974
rect 30156 12870 30212 12908
rect 30380 12964 30436 12974
rect 29596 12796 29764 12852
rect 29484 12350 29486 12402
rect 29538 12350 29540 12402
rect 29484 12338 29540 12350
rect 29596 12180 29652 12190
rect 29372 12124 29540 12180
rect 29372 11956 29428 11966
rect 29260 11954 29428 11956
rect 29260 11902 29374 11954
rect 29426 11902 29428 11954
rect 29260 11900 29428 11902
rect 29260 10500 29316 11900
rect 29372 11890 29428 11900
rect 29484 11284 29540 12124
rect 29596 12086 29652 12124
rect 29708 11732 29764 12796
rect 29932 12850 30100 12852
rect 29932 12798 29934 12850
rect 29986 12798 30100 12850
rect 29932 12796 30100 12798
rect 29932 12786 29988 12796
rect 29932 12628 29988 12638
rect 29820 12404 29876 12414
rect 29820 12290 29876 12348
rect 29820 12238 29822 12290
rect 29874 12238 29876 12290
rect 29820 12226 29876 12238
rect 29708 11666 29764 11676
rect 29596 11284 29652 11294
rect 29484 11282 29652 11284
rect 29484 11230 29598 11282
rect 29650 11230 29652 11282
rect 29484 11228 29652 11230
rect 29036 9102 29038 9154
rect 29090 9102 29092 9154
rect 29036 9090 29092 9102
rect 29148 10498 29316 10500
rect 29148 10446 29262 10498
rect 29314 10446 29316 10498
rect 29148 10444 29316 10446
rect 29036 8596 29092 8606
rect 29036 7474 29092 8540
rect 29036 7422 29038 7474
rect 29090 7422 29092 7474
rect 29036 6132 29092 7422
rect 29036 4676 29092 6076
rect 29148 5348 29204 10444
rect 29260 10434 29316 10444
rect 29596 10052 29652 11228
rect 29820 11172 29876 11182
rect 29372 9828 29428 9838
rect 29260 9268 29316 9278
rect 29260 7140 29316 9212
rect 29372 8148 29428 9772
rect 29596 9828 29652 9996
rect 29596 9762 29652 9772
rect 29708 10948 29764 10958
rect 29484 9602 29540 9614
rect 29484 9550 29486 9602
rect 29538 9550 29540 9602
rect 29484 8596 29540 9550
rect 29596 9268 29652 9278
rect 29596 9154 29652 9212
rect 29708 9266 29764 10892
rect 29820 10834 29876 11116
rect 29820 10782 29822 10834
rect 29874 10782 29876 10834
rect 29820 10770 29876 10782
rect 29708 9214 29710 9266
rect 29762 9214 29764 9266
rect 29708 9202 29764 9214
rect 29820 10164 29876 10174
rect 29596 9102 29598 9154
rect 29650 9102 29652 9154
rect 29596 8932 29652 9102
rect 29596 8866 29652 8876
rect 29484 8530 29540 8540
rect 29596 8372 29652 8382
rect 29820 8372 29876 10108
rect 29932 9042 29988 12572
rect 30380 12180 30436 12908
rect 30380 11956 30436 12124
rect 30492 12178 30548 13804
rect 30604 12852 30660 12862
rect 30604 12402 30660 12796
rect 30716 12850 30772 12862
rect 30716 12798 30718 12850
rect 30770 12798 30772 12850
rect 30716 12740 30772 12798
rect 30828 12852 30884 14812
rect 31276 14756 31332 14766
rect 31276 14662 31332 14700
rect 31388 14530 31444 15092
rect 31388 14478 31390 14530
rect 31442 14478 31444 14530
rect 31388 14466 31444 14478
rect 31276 14308 31332 14318
rect 31612 14308 31668 15486
rect 31724 15426 31780 16604
rect 31836 16436 31892 16446
rect 31836 16100 31892 16380
rect 31836 16006 31892 16044
rect 31724 15374 31726 15426
rect 31778 15374 31780 15426
rect 31724 15362 31780 15374
rect 32060 15204 32116 17164
rect 32172 17108 32228 17118
rect 32172 17014 32228 17052
rect 32284 15652 32340 18958
rect 32396 18452 32452 20132
rect 32508 18452 32564 22316
rect 33404 22148 33460 22158
rect 33068 22146 33460 22148
rect 33068 22094 33406 22146
rect 33458 22094 33460 22146
rect 33068 22092 33460 22094
rect 32732 21474 32788 21486
rect 32732 21422 32734 21474
rect 32786 21422 32788 21474
rect 32620 21364 32676 21374
rect 32620 20914 32676 21308
rect 32620 20862 32622 20914
rect 32674 20862 32676 20914
rect 32620 20850 32676 20862
rect 32620 20580 32676 20590
rect 32620 20244 32676 20524
rect 32620 20178 32676 20188
rect 32732 20020 32788 21422
rect 33068 20914 33124 22092
rect 33404 22082 33460 22092
rect 33516 21924 33572 22316
rect 33740 22148 33796 22158
rect 33740 22054 33796 22092
rect 33068 20862 33070 20914
rect 33122 20862 33124 20914
rect 32620 19964 32788 20020
rect 32844 20244 32900 20254
rect 32620 19796 32676 19964
rect 32844 19908 32900 20188
rect 33068 20020 33124 20862
rect 33404 21868 33572 21924
rect 34300 22036 34356 22046
rect 33404 20188 33460 21868
rect 33740 21812 33796 21822
rect 33628 21474 33684 21486
rect 33628 21422 33630 21474
rect 33682 21422 33684 21474
rect 33516 21026 33572 21038
rect 33516 20974 33518 21026
rect 33570 20974 33572 21026
rect 33516 20916 33572 20974
rect 33516 20822 33572 20860
rect 33068 19954 33124 19964
rect 33292 20132 33460 20188
rect 32620 18676 32676 19740
rect 32620 18610 32676 18620
rect 32732 19906 32900 19908
rect 32732 19854 32846 19906
rect 32898 19854 32900 19906
rect 32732 19852 32900 19854
rect 32508 18396 32676 18452
rect 32396 18340 32452 18396
rect 32396 18338 32564 18340
rect 32396 18286 32398 18338
rect 32450 18286 32564 18338
rect 32396 18284 32564 18286
rect 32396 18274 32452 18284
rect 32508 17668 32564 18284
rect 32508 17574 32564 17612
rect 32620 17220 32676 18396
rect 32732 18340 32788 19852
rect 32844 19842 32900 19852
rect 33292 19236 33348 20132
rect 33516 20020 33572 20030
rect 33516 19926 33572 19964
rect 33628 19908 33684 21422
rect 33628 19684 33684 19852
rect 33180 19180 33348 19236
rect 33516 19628 33684 19684
rect 33516 19236 33572 19628
rect 33740 19460 33796 21756
rect 34300 21812 34356 21980
rect 34524 22036 34580 22990
rect 34860 23042 34916 23054
rect 34860 22990 34862 23042
rect 34914 22990 34916 23042
rect 34524 21970 34580 21980
rect 34748 22146 34804 22158
rect 34748 22094 34750 22146
rect 34802 22094 34804 22146
rect 34300 21746 34356 21756
rect 34076 21588 34132 21598
rect 34076 21494 34132 21532
rect 34412 21476 34468 21486
rect 34300 21474 34468 21476
rect 34300 21422 34414 21474
rect 34466 21422 34468 21474
rect 34300 21420 34468 21422
rect 34300 20916 34356 21420
rect 34412 21410 34468 21420
rect 33964 20580 34020 20590
rect 33964 20486 34020 20524
rect 34300 20580 34356 20860
rect 34412 21026 34468 21038
rect 34412 20974 34414 21026
rect 34466 20974 34468 21026
rect 34412 20914 34468 20974
rect 34412 20862 34414 20914
rect 34466 20862 34468 20914
rect 34412 20850 34468 20862
rect 34300 20514 34356 20524
rect 34412 20020 34468 20030
rect 34300 19964 34412 20020
rect 33964 19908 34020 19918
rect 33964 19814 34020 19852
rect 33628 19348 33684 19358
rect 33740 19348 33796 19404
rect 33628 19346 33796 19348
rect 33628 19294 33630 19346
rect 33682 19294 33796 19346
rect 33628 19292 33796 19294
rect 33628 19282 33684 19292
rect 32732 18274 32788 18284
rect 32844 19012 32900 19022
rect 32620 17154 32676 17164
rect 32396 16996 32452 17006
rect 32396 16902 32452 16940
rect 32508 16882 32564 16894
rect 32508 16830 32510 16882
rect 32562 16830 32564 16882
rect 32508 16100 32564 16830
rect 32508 16034 32564 16044
rect 32732 16884 32788 16894
rect 32284 15586 32340 15596
rect 32620 15986 32676 15998
rect 32620 15934 32622 15986
rect 32674 15934 32676 15986
rect 32620 15652 32676 15934
rect 32620 15586 32676 15596
rect 31276 14306 31668 14308
rect 31276 14254 31278 14306
rect 31330 14254 31668 14306
rect 31276 14252 31668 14254
rect 31948 15148 32116 15204
rect 32172 15428 32228 15438
rect 32172 15148 32228 15372
rect 32396 15428 32452 15438
rect 32396 15426 32564 15428
rect 32396 15374 32398 15426
rect 32450 15374 32564 15426
rect 32396 15372 32564 15374
rect 32396 15362 32452 15372
rect 32284 15316 32340 15326
rect 32284 15222 32340 15260
rect 32508 15316 32564 15372
rect 32508 15250 32564 15260
rect 32396 15204 32452 15214
rect 31276 14242 31332 14252
rect 31052 13076 31108 13086
rect 31052 12962 31108 13020
rect 31052 12910 31054 12962
rect 31106 12910 31108 12962
rect 31052 12898 31108 12910
rect 30828 12850 30996 12852
rect 30828 12798 30830 12850
rect 30882 12798 30996 12850
rect 30828 12796 30996 12798
rect 30828 12786 30884 12796
rect 30716 12674 30772 12684
rect 30604 12350 30606 12402
rect 30658 12350 30660 12402
rect 30604 12338 30660 12350
rect 30716 12516 30772 12526
rect 30492 12126 30494 12178
rect 30546 12126 30548 12178
rect 30492 12114 30548 12126
rect 30716 12066 30772 12460
rect 30940 12516 30996 12796
rect 31500 12850 31556 12862
rect 31500 12798 31502 12850
rect 31554 12798 31556 12850
rect 31500 12740 31556 12798
rect 31612 12852 31668 12862
rect 31612 12758 31668 12796
rect 31836 12740 31892 12750
rect 31500 12674 31556 12684
rect 31724 12738 31892 12740
rect 31724 12686 31838 12738
rect 31890 12686 31892 12738
rect 31724 12684 31892 12686
rect 30940 12450 30996 12460
rect 31612 12404 31668 12414
rect 30940 12180 30996 12218
rect 30940 12114 30996 12124
rect 30716 12014 30718 12066
rect 30770 12014 30772 12066
rect 30716 12002 30772 12014
rect 30828 12068 30884 12078
rect 30156 11900 30436 11956
rect 30044 11732 30100 11742
rect 30044 11170 30100 11676
rect 30156 11396 30212 11900
rect 30604 11788 30660 11798
rect 30156 11394 30548 11396
rect 30156 11342 30158 11394
rect 30210 11342 30548 11394
rect 30156 11340 30548 11342
rect 30156 11330 30212 11340
rect 30044 11118 30046 11170
rect 30098 11118 30100 11170
rect 30044 11060 30100 11118
rect 30044 10994 30100 11004
rect 30492 10834 30548 11340
rect 30492 10782 30494 10834
rect 30546 10782 30548 10834
rect 30492 10770 30548 10782
rect 30604 10610 30660 11732
rect 30828 11396 30884 12012
rect 31052 12068 31108 12078
rect 31052 11956 31108 12012
rect 31500 12068 31556 12078
rect 30604 10558 30606 10610
rect 30658 10558 30660 10610
rect 30604 10546 30660 10558
rect 30716 11340 30884 11396
rect 30940 11900 31108 11956
rect 31164 11956 31220 11994
rect 30716 10164 30772 11340
rect 30828 11172 30884 11182
rect 30828 11078 30884 11116
rect 30492 10108 30772 10164
rect 30268 10052 30324 10062
rect 30268 9958 30324 9996
rect 30044 9940 30100 9950
rect 30044 9846 30100 9884
rect 29932 8990 29934 9042
rect 29986 8990 29988 9042
rect 29932 8978 29988 8990
rect 30156 9604 30212 9614
rect 29596 8278 29652 8316
rect 29708 8370 29876 8372
rect 29708 8318 29822 8370
rect 29874 8318 29876 8370
rect 29708 8316 29876 8318
rect 29372 8092 29652 8148
rect 29260 7074 29316 7084
rect 29372 7700 29428 7710
rect 29260 6020 29316 6030
rect 29260 5926 29316 5964
rect 29148 5282 29204 5292
rect 29372 5684 29428 7644
rect 29596 7476 29652 8092
rect 29708 8036 29764 8316
rect 29820 8306 29876 8316
rect 29708 7970 29764 7980
rect 29820 8034 29876 8046
rect 29820 7982 29822 8034
rect 29874 7982 29876 8034
rect 29708 7700 29764 7710
rect 29708 7606 29764 7644
rect 29596 7362 29652 7420
rect 29596 7310 29598 7362
rect 29650 7310 29652 7362
rect 29596 7298 29652 7310
rect 29820 6916 29876 7982
rect 29820 6850 29876 6860
rect 29932 7250 29988 7262
rect 29932 7198 29934 7250
rect 29986 7198 29988 7250
rect 29932 7028 29988 7198
rect 29932 6804 29988 6972
rect 29932 6738 29988 6748
rect 30156 6690 30212 9548
rect 30492 8372 30548 10108
rect 30604 9940 30660 9950
rect 30604 9846 30660 9884
rect 30828 9716 30884 9726
rect 30828 9154 30884 9660
rect 30828 9102 30830 9154
rect 30882 9102 30884 9154
rect 30828 9090 30884 9102
rect 30492 7700 30548 8316
rect 30604 8036 30660 8074
rect 30604 7970 30660 7980
rect 30940 7924 30996 11900
rect 31164 11890 31220 11900
rect 31164 11788 31220 11798
rect 31220 11732 31332 11788
rect 31500 11732 31556 12012
rect 31164 11722 31220 11732
rect 31276 11676 31556 11732
rect 31164 11396 31220 11406
rect 31164 10834 31220 11340
rect 31388 11282 31444 11294
rect 31388 11230 31390 11282
rect 31442 11230 31444 11282
rect 31388 10948 31444 11230
rect 31388 10882 31444 10892
rect 31164 10782 31166 10834
rect 31218 10782 31220 10834
rect 31164 10770 31220 10782
rect 31388 10724 31444 10734
rect 31388 10630 31444 10668
rect 31500 10612 31556 10622
rect 31500 10518 31556 10556
rect 31388 10276 31444 10286
rect 31164 9940 31220 9950
rect 31164 9714 31220 9884
rect 31164 9662 31166 9714
rect 31218 9662 31220 9714
rect 31164 9650 31220 9662
rect 31388 9826 31444 10220
rect 31612 10052 31668 12348
rect 31388 9774 31390 9826
rect 31442 9774 31444 9826
rect 31052 9604 31108 9614
rect 31052 9510 31108 9548
rect 31276 9604 31332 9614
rect 31276 9492 31332 9548
rect 31164 9436 31332 9492
rect 31052 9268 31108 9278
rect 31164 9268 31220 9436
rect 31052 9266 31220 9268
rect 31052 9214 31054 9266
rect 31106 9214 31220 9266
rect 31052 9212 31220 9214
rect 31276 9268 31332 9278
rect 31388 9268 31444 9774
rect 31276 9266 31444 9268
rect 31276 9214 31278 9266
rect 31330 9214 31444 9266
rect 31276 9212 31444 9214
rect 31500 9996 31668 10052
rect 31052 9202 31108 9212
rect 31276 9202 31332 9212
rect 30940 7858 30996 7868
rect 31164 9044 31220 9054
rect 30492 7634 30548 7644
rect 30604 7812 30660 7822
rect 30604 7698 30660 7756
rect 30604 7646 30606 7698
rect 30658 7646 30660 7698
rect 30492 7476 30548 7486
rect 30492 7382 30548 7420
rect 30604 7364 30660 7646
rect 30828 7476 30884 7514
rect 30828 7410 30884 7420
rect 31164 7364 31220 8988
rect 31388 9044 31444 9054
rect 31388 8950 31444 8988
rect 31500 8596 31556 9996
rect 31612 9828 31668 9838
rect 31612 9734 31668 9772
rect 31724 9268 31780 12684
rect 31836 12674 31892 12684
rect 31948 12628 32004 15148
rect 32172 15092 32340 15148
rect 32172 14980 32228 14990
rect 32060 14420 32116 14430
rect 32060 13636 32116 14364
rect 32172 14418 32228 14924
rect 32284 14532 32340 15092
rect 32396 15090 32452 15148
rect 32396 15038 32398 15090
rect 32450 15038 32452 15090
rect 32396 15026 32452 15038
rect 32732 14642 32788 16828
rect 32844 16660 32900 18956
rect 32844 16594 32900 16604
rect 32956 18340 33012 18350
rect 32844 16100 32900 16110
rect 32844 15652 32900 16044
rect 32956 15988 33012 18284
rect 33180 17780 33236 19180
rect 33516 19170 33572 19180
rect 34188 19236 34244 19246
rect 34188 19142 34244 19180
rect 33292 19012 33348 19022
rect 33292 18918 33348 18956
rect 33516 18340 33572 18350
rect 34076 18340 34132 18378
rect 33516 18338 33684 18340
rect 33516 18286 33518 18338
rect 33570 18286 33684 18338
rect 33516 18284 33684 18286
rect 33516 18274 33572 18284
rect 33180 17724 33348 17780
rect 33180 17554 33236 17566
rect 33180 17502 33182 17554
rect 33234 17502 33236 17554
rect 33068 17444 33124 17454
rect 33068 16098 33124 17388
rect 33180 16210 33236 17502
rect 33292 16548 33348 17724
rect 33628 17668 33684 18284
rect 34076 18274 34132 18284
rect 33628 16882 33684 17612
rect 34076 18116 34132 18126
rect 33628 16830 33630 16882
rect 33682 16830 33684 16882
rect 33628 16818 33684 16830
rect 33740 16996 33796 17006
rect 33292 16482 33348 16492
rect 33180 16158 33182 16210
rect 33234 16158 33236 16210
rect 33180 16146 33236 16158
rect 33404 16212 33460 16222
rect 33068 16046 33070 16098
rect 33122 16046 33124 16098
rect 33068 16034 33124 16046
rect 33292 16100 33348 16110
rect 33404 16100 33460 16156
rect 33292 16098 33460 16100
rect 33292 16046 33294 16098
rect 33346 16046 33460 16098
rect 33292 16044 33460 16046
rect 33628 16212 33684 16222
rect 33292 16034 33348 16044
rect 32956 15876 33012 15932
rect 32956 15820 33236 15876
rect 32844 15586 32900 15596
rect 32732 14590 32734 14642
rect 32786 14590 32788 14642
rect 32732 14578 32788 14590
rect 32396 14532 32452 14542
rect 32620 14532 32676 14542
rect 32284 14530 32564 14532
rect 32284 14478 32398 14530
rect 32450 14478 32564 14530
rect 32284 14476 32564 14478
rect 32396 14466 32452 14476
rect 32172 14366 32174 14418
rect 32226 14366 32228 14418
rect 32172 14084 32228 14366
rect 32508 14084 32564 14476
rect 32620 14438 32676 14476
rect 32844 14532 32900 14542
rect 32844 14530 33012 14532
rect 32844 14478 32846 14530
rect 32898 14478 33012 14530
rect 32844 14476 33012 14478
rect 32844 14466 32900 14476
rect 32228 14028 32340 14084
rect 32508 14028 32788 14084
rect 32172 14018 32228 14028
rect 32060 13504 32116 13580
rect 31948 12562 32004 12572
rect 32060 13076 32116 13086
rect 32060 12404 32116 13020
rect 31948 12348 32116 12404
rect 31836 12178 31892 12190
rect 31836 12126 31838 12178
rect 31890 12126 31892 12178
rect 31836 10948 31892 12126
rect 31836 10882 31892 10892
rect 31948 11282 32004 12348
rect 32284 12068 32340 14028
rect 32732 13970 32788 14028
rect 32732 13918 32734 13970
rect 32786 13918 32788 13970
rect 32732 13906 32788 13918
rect 32844 13972 32900 13982
rect 32508 13860 32564 13870
rect 32508 13766 32564 13804
rect 32844 13858 32900 13916
rect 32844 13806 32846 13858
rect 32898 13806 32900 13858
rect 32844 13794 32900 13806
rect 32732 13748 32788 13758
rect 32396 13524 32452 13534
rect 32396 12962 32452 13468
rect 32396 12910 32398 12962
rect 32450 12910 32452 12962
rect 32396 12898 32452 12910
rect 32732 12404 32788 13692
rect 32844 12404 32900 12414
rect 32732 12402 32900 12404
rect 32732 12350 32846 12402
rect 32898 12350 32900 12402
rect 32732 12348 32900 12350
rect 32844 12338 32900 12348
rect 31948 11230 31950 11282
rect 32002 11230 32004 11282
rect 31948 9604 32004 11230
rect 32060 12066 32340 12068
rect 32060 12014 32286 12066
rect 32338 12014 32340 12066
rect 32060 12012 32340 12014
rect 32060 10722 32116 12012
rect 32284 12002 32340 12012
rect 32956 11732 33012 14476
rect 33068 13412 33124 13422
rect 33068 13074 33124 13356
rect 33068 13022 33070 13074
rect 33122 13022 33124 13074
rect 33068 13010 33124 13022
rect 32956 11666 33012 11676
rect 33068 12292 33124 12302
rect 32060 10670 32062 10722
rect 32114 10670 32116 10722
rect 32060 10658 32116 10670
rect 32172 11506 32228 11518
rect 32172 11454 32174 11506
rect 32226 11454 32228 11506
rect 31948 9538 32004 9548
rect 32060 9492 32116 9502
rect 31836 9268 31892 9278
rect 31724 9266 31892 9268
rect 31724 9214 31838 9266
rect 31890 9214 31892 9266
rect 31724 9212 31892 9214
rect 31836 9202 31892 9212
rect 32060 9266 32116 9436
rect 32060 9214 32062 9266
rect 32114 9214 32116 9266
rect 31724 8820 31780 8830
rect 31276 8540 31556 8596
rect 31612 8818 31780 8820
rect 31612 8766 31726 8818
rect 31778 8766 31780 8818
rect 31612 8764 31780 8766
rect 31276 7812 31332 8540
rect 31388 8372 31444 8382
rect 31388 8278 31444 8316
rect 31612 8260 31668 8764
rect 31724 8754 31780 8764
rect 31724 8596 31780 8606
rect 31724 8370 31780 8540
rect 32060 8484 32116 9214
rect 32172 9268 32228 11454
rect 32732 11508 32788 11518
rect 32284 11060 32340 11070
rect 32732 11060 32788 11452
rect 32844 11396 32900 11406
rect 32844 11302 32900 11340
rect 32956 11284 33012 11294
rect 33068 11284 33124 12236
rect 33180 11396 33236 15820
rect 33516 15316 33572 15326
rect 33516 15222 33572 15260
rect 33628 15148 33684 16156
rect 33740 15652 33796 16940
rect 33852 16436 33908 16446
rect 33852 16322 33908 16380
rect 33852 16270 33854 16322
rect 33906 16270 33908 16322
rect 33852 16258 33908 16270
rect 33964 15986 34020 15998
rect 33964 15934 33966 15986
rect 34018 15934 34020 15986
rect 33740 15596 33908 15652
rect 33740 15426 33796 15438
rect 33740 15374 33742 15426
rect 33794 15374 33796 15426
rect 33740 15316 33796 15374
rect 33740 15250 33796 15260
rect 33852 15426 33908 15596
rect 33852 15374 33854 15426
rect 33906 15374 33908 15426
rect 33628 15092 33796 15148
rect 33516 14756 33572 14766
rect 33292 14644 33348 14654
rect 33292 14530 33348 14588
rect 33292 14478 33294 14530
rect 33346 14478 33348 14530
rect 33292 14466 33348 14478
rect 33516 14418 33572 14700
rect 33628 14644 33684 14654
rect 33628 14530 33684 14588
rect 33628 14478 33630 14530
rect 33682 14478 33684 14530
rect 33628 14466 33684 14478
rect 33516 14366 33518 14418
rect 33570 14366 33572 14418
rect 33180 11330 33236 11340
rect 33292 13748 33348 13758
rect 32956 11282 33124 11284
rect 32956 11230 32958 11282
rect 33010 11230 33124 11282
rect 32956 11228 33124 11230
rect 32956 11218 33012 11228
rect 33180 11170 33236 11182
rect 33180 11118 33182 11170
rect 33234 11118 33236 11170
rect 33180 11060 33236 11118
rect 32732 11004 33236 11060
rect 32284 10834 32340 11004
rect 32284 10782 32286 10834
rect 32338 10782 32340 10834
rect 32284 10770 32340 10782
rect 32620 10836 32676 10846
rect 32620 10742 32676 10780
rect 32508 10610 32564 10622
rect 32508 10558 32510 10610
rect 32562 10558 32564 10610
rect 32508 10500 32564 10558
rect 32508 10434 32564 10444
rect 32620 10556 33236 10612
rect 32620 10498 32676 10556
rect 32620 10446 32622 10498
rect 32674 10446 32676 10498
rect 32620 10434 32676 10446
rect 32732 10388 32788 10398
rect 32172 9202 32228 9212
rect 32508 9826 32564 9838
rect 32508 9774 32510 9826
rect 32562 9774 32564 9826
rect 32284 9044 32340 9054
rect 32284 8950 32340 8988
rect 32060 8418 32116 8428
rect 31724 8318 31726 8370
rect 31778 8318 31780 8370
rect 31724 8306 31780 8318
rect 31276 7746 31332 7756
rect 31500 8204 31668 8260
rect 32508 8260 32564 9774
rect 32732 9266 32788 10332
rect 33180 9938 33236 10556
rect 33292 10388 33348 13692
rect 33516 13076 33572 14366
rect 33628 14084 33684 14094
rect 33628 13858 33684 14028
rect 33628 13806 33630 13858
rect 33682 13806 33684 13858
rect 33628 13794 33684 13806
rect 33516 13010 33572 13020
rect 33628 13636 33684 13646
rect 33628 12290 33684 13580
rect 33740 12402 33796 15092
rect 33852 14868 33908 15374
rect 33964 15204 34020 15934
rect 34076 15316 34132 18060
rect 34076 15250 34132 15260
rect 34300 15204 34356 19964
rect 34412 19926 34468 19964
rect 34524 19236 34580 19246
rect 34524 18900 34580 19180
rect 34412 16884 34468 16894
rect 34412 16790 34468 16828
rect 34524 15988 34580 18844
rect 34636 19010 34692 19022
rect 34636 18958 34638 19010
rect 34690 18958 34692 19010
rect 34636 17332 34692 18958
rect 34636 17266 34692 17276
rect 34748 17220 34804 22094
rect 34860 21812 34916 22990
rect 35084 22482 35140 23100
rect 35420 23044 35476 23054
rect 35420 23042 35700 23044
rect 35420 22990 35422 23042
rect 35474 22990 35700 23042
rect 35420 22988 35700 22990
rect 35420 22978 35476 22988
rect 35644 22930 35700 22988
rect 35644 22878 35646 22930
rect 35698 22878 35700 22930
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22430 35086 22482
rect 35138 22430 35140 22482
rect 35084 22372 35140 22430
rect 35084 22306 35140 22316
rect 35532 22148 35588 22158
rect 35532 22054 35588 22092
rect 35084 22036 35140 22046
rect 34860 21810 35028 21812
rect 34860 21758 34862 21810
rect 34914 21758 35028 21810
rect 34860 21756 35028 21758
rect 34860 21746 34916 21756
rect 34860 21026 34916 21038
rect 34860 20974 34862 21026
rect 34914 20974 34916 21026
rect 34860 20914 34916 20974
rect 34860 20862 34862 20914
rect 34914 20862 34916 20914
rect 34860 20850 34916 20862
rect 34860 20356 34916 20366
rect 34860 20242 34916 20300
rect 34860 20190 34862 20242
rect 34914 20190 34916 20242
rect 34860 20178 34916 20190
rect 34972 20188 35028 21756
rect 35084 21026 35140 21980
rect 35420 21476 35476 21486
rect 35420 21474 35588 21476
rect 35420 21422 35422 21474
rect 35474 21422 35588 21474
rect 35420 21420 35588 21422
rect 35420 21410 35476 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20974 35086 21026
rect 35138 20974 35140 21026
rect 35084 20962 35140 20974
rect 35308 21026 35364 21038
rect 35308 20974 35310 21026
rect 35362 20974 35364 21026
rect 35308 20914 35364 20974
rect 35308 20862 35310 20914
rect 35362 20862 35364 20914
rect 35308 20188 35364 20862
rect 35532 20580 35588 21420
rect 35644 20916 35700 22878
rect 35868 23042 35924 23054
rect 35868 22990 35870 23042
rect 35922 22990 35924 23042
rect 35868 22036 35924 22990
rect 35980 22594 36036 24556
rect 35980 22542 35982 22594
rect 36034 22542 36036 22594
rect 35980 22530 36036 22542
rect 36204 23042 36260 23054
rect 36204 22990 36206 23042
rect 36258 22990 36260 23042
rect 35868 21970 35924 21980
rect 35980 22146 36036 22158
rect 35980 22094 35982 22146
rect 36034 22094 36036 22146
rect 35756 21924 35812 21934
rect 35756 21812 35812 21868
rect 35756 21810 35924 21812
rect 35756 21758 35758 21810
rect 35810 21758 35924 21810
rect 35756 21756 35924 21758
rect 35756 21746 35812 21756
rect 35756 20916 35812 20926
rect 35644 20860 35756 20916
rect 35756 20822 35812 20860
rect 35532 20514 35588 20524
rect 35868 20580 35924 21756
rect 34972 20132 35812 20188
rect 34972 20020 35028 20132
rect 34972 19954 35028 19964
rect 35084 19908 35140 19918
rect 35084 19346 35140 19852
rect 35420 19908 35476 19918
rect 35420 19906 35588 19908
rect 35420 19854 35422 19906
rect 35474 19854 35588 19906
rect 35420 19852 35588 19854
rect 35420 19842 35476 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 19294 35086 19346
rect 35138 19294 35140 19346
rect 34860 18340 34916 18350
rect 34860 18246 34916 18284
rect 34972 18228 35028 18238
rect 34972 18134 35028 18172
rect 34748 17154 34804 17164
rect 34972 16212 35028 16222
rect 34636 15988 34692 15998
rect 34524 15986 34692 15988
rect 34524 15934 34638 15986
rect 34690 15934 34692 15986
rect 34524 15932 34692 15934
rect 34412 15876 34468 15886
rect 34412 15782 34468 15820
rect 34300 15148 34468 15204
rect 33964 15138 34020 15148
rect 33852 14812 34244 14868
rect 34188 14754 34244 14812
rect 34188 14702 34190 14754
rect 34242 14702 34244 14754
rect 34188 14690 34244 14702
rect 34300 14420 34356 14430
rect 34300 14326 34356 14364
rect 33852 13972 33908 13982
rect 33852 13878 33908 13916
rect 34076 13748 34132 13758
rect 34300 13748 34356 13758
rect 34076 13746 34244 13748
rect 34076 13694 34078 13746
rect 34130 13694 34244 13746
rect 34076 13692 34244 13694
rect 34076 13682 34132 13692
rect 33964 13634 34020 13646
rect 33964 13582 33966 13634
rect 34018 13582 34020 13634
rect 33964 13412 34020 13582
rect 33964 13346 34020 13356
rect 33740 12350 33742 12402
rect 33794 12350 33796 12402
rect 33740 12338 33796 12350
rect 33852 13300 33908 13310
rect 33628 12238 33630 12290
rect 33682 12238 33684 12290
rect 33628 12226 33684 12238
rect 33852 12180 33908 13244
rect 33852 12048 33908 12124
rect 33964 13076 34020 13086
rect 33740 11620 33796 11630
rect 33292 10322 33348 10332
rect 33516 11284 33572 11294
rect 33516 11170 33572 11228
rect 33516 11118 33518 11170
rect 33570 11118 33572 11170
rect 33180 9886 33182 9938
rect 33234 9886 33236 9938
rect 33180 9874 33236 9886
rect 33516 9492 33572 11118
rect 33740 10724 33796 11564
rect 33740 10630 33796 10668
rect 33628 10612 33684 10622
rect 33964 10612 34020 13020
rect 34076 11954 34132 11966
rect 34076 11902 34078 11954
rect 34130 11902 34132 11954
rect 34076 10948 34132 11902
rect 34188 11956 34244 13692
rect 34300 13654 34356 13692
rect 34412 13300 34468 15148
rect 34524 14420 34580 15932
rect 34636 15922 34692 15932
rect 34748 15988 34804 15998
rect 34748 15894 34804 15932
rect 34524 14354 34580 14364
rect 34636 15540 34692 15550
rect 34636 14308 34692 15484
rect 34860 15316 34916 15326
rect 34860 15202 34916 15260
rect 34972 15314 35028 16156
rect 34972 15262 34974 15314
rect 35026 15262 35028 15314
rect 34972 15250 35028 15262
rect 34860 15150 34862 15202
rect 34914 15150 34916 15202
rect 34860 15138 34916 15150
rect 34860 14868 34916 14878
rect 34860 14644 34916 14812
rect 35084 14644 35140 19294
rect 35532 19236 35588 19852
rect 35756 19906 35812 20132
rect 35756 19854 35758 19906
rect 35810 19854 35812 19906
rect 35756 19572 35812 19854
rect 35756 19506 35812 19516
rect 35420 18340 35476 18350
rect 35420 18246 35476 18284
rect 35532 18226 35588 19180
rect 35756 19012 35812 19022
rect 35532 18174 35534 18226
rect 35586 18174 35588 18226
rect 35532 18162 35588 18174
rect 35644 18956 35756 19012
rect 35644 18788 35700 18956
rect 35756 18918 35812 18956
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35308 17780 35364 17790
rect 35308 17778 35588 17780
rect 35308 17726 35310 17778
rect 35362 17726 35588 17778
rect 35308 17724 35588 17726
rect 35308 17714 35364 17724
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16212 35364 16222
rect 35308 16098 35364 16156
rect 35308 16046 35310 16098
rect 35362 16046 35364 16098
rect 35308 16034 35364 16046
rect 35420 15988 35476 15998
rect 35532 15988 35588 17724
rect 35644 16660 35700 18732
rect 35868 18564 35924 20524
rect 35868 18498 35924 18508
rect 35868 18338 35924 18350
rect 35868 18286 35870 18338
rect 35922 18286 35924 18338
rect 35868 18226 35924 18286
rect 35868 18174 35870 18226
rect 35922 18174 35924 18226
rect 35868 18162 35924 18174
rect 35980 18228 36036 22094
rect 36204 21026 36260 22990
rect 36316 22260 36372 27020
rect 43260 25284 43316 25294
rect 38444 24836 38500 24846
rect 36876 24052 36932 24062
rect 36876 23958 36932 23996
rect 37548 24052 37604 24062
rect 36428 23716 36484 23726
rect 36428 23714 36708 23716
rect 36428 23662 36430 23714
rect 36482 23662 36708 23714
rect 36428 23660 36708 23662
rect 36428 23650 36484 23660
rect 36428 22708 36484 22718
rect 36428 22594 36484 22652
rect 36428 22542 36430 22594
rect 36482 22542 36484 22594
rect 36428 22482 36484 22542
rect 36428 22430 36430 22482
rect 36482 22430 36484 22482
rect 36428 22418 36484 22430
rect 36540 22596 36596 22606
rect 36316 22204 36484 22260
rect 36204 20974 36206 21026
rect 36258 20974 36260 21026
rect 36204 20962 36260 20974
rect 36316 21474 36372 21486
rect 36316 21422 36318 21474
rect 36370 21422 36372 21474
rect 36092 20916 36148 20926
rect 36092 20804 36148 20860
rect 36204 20804 36260 20814
rect 36092 20802 36260 20804
rect 36092 20750 36206 20802
rect 36258 20750 36260 20802
rect 36092 20748 36260 20750
rect 36204 20738 36260 20748
rect 36204 20468 36260 20478
rect 36204 20188 36260 20412
rect 36316 20356 36372 21422
rect 36316 20290 36372 20300
rect 36204 20132 36372 20188
rect 36204 19906 36260 19918
rect 36204 19854 36206 19906
rect 36258 19854 36260 19906
rect 36204 19796 36260 19854
rect 36204 19730 36260 19740
rect 36204 19010 36260 19022
rect 36204 18958 36206 19010
rect 36258 18958 36260 19010
rect 35980 18162 36036 18172
rect 36092 18450 36148 18462
rect 36092 18398 36094 18450
rect 36146 18398 36148 18450
rect 36092 17668 36148 18398
rect 35980 17612 36148 17668
rect 35980 17554 36036 17612
rect 35980 17502 35982 17554
rect 36034 17502 36036 17554
rect 35644 16604 35924 16660
rect 35476 15932 35588 15988
rect 35644 16436 35700 16446
rect 35644 16098 35700 16380
rect 35644 16046 35646 16098
rect 35698 16046 35700 16098
rect 35420 15894 35476 15932
rect 35644 15764 35700 16046
rect 35644 15698 35700 15708
rect 35756 16212 35812 16222
rect 35644 15540 35700 15550
rect 35644 15446 35700 15484
rect 35532 15316 35588 15326
rect 35532 15222 35588 15260
rect 35644 15204 35700 15214
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34860 14642 35140 14644
rect 34860 14590 34862 14642
rect 34914 14590 35140 14642
rect 34860 14588 35140 14590
rect 34860 14578 34916 14588
rect 34636 14252 34916 14308
rect 34860 13970 34916 14252
rect 34972 14306 35028 14318
rect 34972 14254 34974 14306
rect 35026 14254 35028 14306
rect 34972 14196 35028 14254
rect 34972 14130 35028 14140
rect 35420 14306 35476 14318
rect 35420 14254 35422 14306
rect 35474 14254 35476 14306
rect 34860 13918 34862 13970
rect 34914 13918 34916 13970
rect 34860 13906 34916 13918
rect 34748 13636 34804 13646
rect 34412 13244 34692 13300
rect 34188 11890 34244 11900
rect 34300 12292 34356 12302
rect 34188 11284 34244 11294
rect 34300 11284 34356 12236
rect 34524 12292 34580 12302
rect 34524 12198 34580 12236
rect 34412 11844 34468 11854
rect 34412 11508 34468 11788
rect 34412 11442 34468 11452
rect 34524 11732 34580 11742
rect 34412 11284 34468 11294
rect 34300 11282 34468 11284
rect 34300 11230 34414 11282
rect 34466 11230 34468 11282
rect 34300 11228 34468 11230
rect 34188 11190 34244 11228
rect 34412 10948 34468 11228
rect 34524 11170 34580 11676
rect 34524 11118 34526 11170
rect 34578 11118 34580 11170
rect 34524 11106 34580 11118
rect 34636 11394 34692 13244
rect 34636 11342 34638 11394
rect 34690 11342 34692 11394
rect 34636 10948 34692 11342
rect 34412 10892 34580 10948
rect 34076 10882 34132 10892
rect 34300 10836 34356 10846
rect 34300 10742 34356 10780
rect 34412 10612 34468 10622
rect 33964 10610 34468 10612
rect 33964 10558 34414 10610
rect 34466 10558 34468 10610
rect 33964 10556 34468 10558
rect 33628 10518 33684 10556
rect 34412 10546 34468 10556
rect 34524 10612 34580 10892
rect 34636 10882 34692 10892
rect 33516 9426 33572 9436
rect 33740 10386 33796 10398
rect 33740 10334 33742 10386
rect 33794 10334 33796 10386
rect 33740 9380 33796 10334
rect 34300 10164 34356 10174
rect 33740 9314 33796 9324
rect 33964 10052 34020 10062
rect 32732 9214 32734 9266
rect 32786 9214 32788 9266
rect 32732 9202 32788 9214
rect 33852 9268 33908 9278
rect 33852 9174 33908 9212
rect 33964 8930 34020 9996
rect 33964 8878 33966 8930
rect 34018 8878 34020 8930
rect 33964 8866 34020 8878
rect 33628 8818 33684 8830
rect 33628 8766 33630 8818
rect 33682 8766 33684 8818
rect 33628 8596 33684 8766
rect 33628 8530 33684 8540
rect 33404 8372 33460 8382
rect 33404 8278 33460 8316
rect 32620 8260 32676 8270
rect 32508 8258 32676 8260
rect 32508 8206 32622 8258
rect 32674 8206 32676 8258
rect 32508 8204 32676 8206
rect 31276 7364 31332 7374
rect 31164 7362 31332 7364
rect 31164 7310 31278 7362
rect 31330 7310 31332 7362
rect 31164 7308 31332 7310
rect 30604 7298 30660 7308
rect 31276 7298 31332 7308
rect 30156 6638 30158 6690
rect 30210 6638 30212 6690
rect 30156 6626 30212 6638
rect 30380 6692 30436 6702
rect 31388 6692 31444 6702
rect 31500 6692 31556 8204
rect 31612 8034 31668 8046
rect 31612 7982 31614 8034
rect 31666 7982 31668 8034
rect 31612 7924 31668 7982
rect 31612 7858 31668 7868
rect 32508 7812 32564 7822
rect 31724 7698 31780 7710
rect 31724 7646 31726 7698
rect 31778 7646 31780 7698
rect 30380 6690 30884 6692
rect 30380 6638 30382 6690
rect 30434 6638 30884 6690
rect 30380 6636 30884 6638
rect 30380 6626 30436 6636
rect 29708 6580 29764 6590
rect 29708 6486 29764 6524
rect 29932 6466 29988 6478
rect 29932 6414 29934 6466
rect 29986 6414 29988 6466
rect 29932 6356 29988 6414
rect 29932 6290 29988 6300
rect 30044 6466 30100 6478
rect 30044 6414 30046 6466
rect 30098 6414 30100 6466
rect 29036 4610 29092 4620
rect 29372 4226 29428 5628
rect 29372 4174 29374 4226
rect 29426 4174 29428 4226
rect 29372 4162 29428 4174
rect 29708 5010 29764 5022
rect 29708 4958 29710 5010
rect 29762 4958 29764 5010
rect 28588 3666 28980 3668
rect 28588 3614 28590 3666
rect 28642 3614 28980 3666
rect 28588 3612 28980 3614
rect 29260 3668 29316 3678
rect 28588 3602 28644 3612
rect 29260 3574 29316 3612
rect 29708 3388 29764 4958
rect 30044 4452 30100 6414
rect 30828 6132 30884 6636
rect 31388 6690 31556 6692
rect 31388 6638 31390 6690
rect 31442 6638 31556 6690
rect 31388 6636 31556 6638
rect 31612 6692 31668 6702
rect 31724 6692 31780 7646
rect 32508 7586 32564 7756
rect 32508 7534 32510 7586
rect 32562 7534 32564 7586
rect 32508 7522 32564 7534
rect 31612 6690 31780 6692
rect 31612 6638 31614 6690
rect 31666 6638 31780 6690
rect 31612 6636 31780 6638
rect 31836 7474 31892 7486
rect 31836 7422 31838 7474
rect 31890 7422 31892 7474
rect 31388 6626 31444 6636
rect 31612 6626 31668 6636
rect 30940 6580 30996 6590
rect 30940 6486 30996 6524
rect 31276 6580 31332 6590
rect 31276 6486 31332 6524
rect 31164 6466 31220 6478
rect 31164 6414 31166 6466
rect 31218 6414 31220 6466
rect 30940 6132 30996 6142
rect 30828 6130 30996 6132
rect 30828 6078 30942 6130
rect 30994 6078 30996 6130
rect 30828 6076 30996 6078
rect 30940 6066 30996 6076
rect 30492 5906 30548 5918
rect 30492 5854 30494 5906
rect 30546 5854 30548 5906
rect 30492 5572 30548 5854
rect 30940 5908 30996 5918
rect 30940 5814 30996 5852
rect 31052 5796 31108 5806
rect 31052 5702 31108 5740
rect 30492 5506 30548 5516
rect 31052 5236 31108 5246
rect 31052 5142 31108 5180
rect 30828 5012 30884 5022
rect 30044 4386 30100 4396
rect 30716 4452 30772 4462
rect 30716 4358 30772 4396
rect 29932 4340 29988 4350
rect 29932 4246 29988 4284
rect 25788 1586 25844 1596
rect 26684 800 26740 3388
rect 28028 3332 28532 3388
rect 29372 3332 29764 3388
rect 30268 3444 30324 3482
rect 30828 3388 30884 4956
rect 30268 3378 30324 3388
rect 30716 3332 30884 3388
rect 28028 800 28084 3332
rect 29372 2660 29428 3332
rect 29372 800 29428 2604
rect 30716 800 30772 3332
rect 31164 2548 31220 6414
rect 31500 5908 31556 5918
rect 31276 5794 31332 5806
rect 31276 5742 31278 5794
rect 31330 5742 31332 5794
rect 31276 5460 31332 5742
rect 31276 5394 31332 5404
rect 31388 5572 31444 5582
rect 31388 3554 31444 5516
rect 31500 5236 31556 5852
rect 31724 5796 31780 5806
rect 31724 5348 31780 5740
rect 31836 5684 31892 7422
rect 32060 7364 32116 7374
rect 31836 5618 31892 5628
rect 31948 7362 32116 7364
rect 31948 7310 32062 7362
rect 32114 7310 32116 7362
rect 31948 7308 32116 7310
rect 31948 5460 32004 7308
rect 32060 7298 32116 7308
rect 32284 7252 32340 7262
rect 32284 7140 32340 7196
rect 32060 7084 32340 7140
rect 32060 5796 32116 7084
rect 32060 5730 32116 5740
rect 32284 6692 32340 6702
rect 32620 6692 32676 8204
rect 33740 8036 33796 8046
rect 33068 7924 33124 7934
rect 32284 6690 32676 6692
rect 32284 6638 32286 6690
rect 32338 6638 32676 6690
rect 32284 6636 32676 6638
rect 32844 7474 32900 7486
rect 32844 7422 32846 7474
rect 32898 7422 32900 7474
rect 32172 5682 32228 5694
rect 32172 5630 32174 5682
rect 32226 5630 32228 5682
rect 32060 5460 32116 5470
rect 31948 5404 32060 5460
rect 31724 5292 32004 5348
rect 31612 5236 31668 5246
rect 31500 5234 31668 5236
rect 31500 5182 31614 5234
rect 31666 5182 31668 5234
rect 31500 5180 31668 5182
rect 31612 5170 31668 5180
rect 31388 3502 31390 3554
rect 31442 3502 31444 3554
rect 31388 3490 31444 3502
rect 31836 4228 31892 4238
rect 31836 3554 31892 4172
rect 31948 3778 32004 5292
rect 31948 3726 31950 3778
rect 32002 3726 32004 3778
rect 31948 3714 32004 3726
rect 32060 3668 32116 5404
rect 32172 5236 32228 5630
rect 32172 5170 32228 5180
rect 32284 4340 32340 6636
rect 32732 6132 32788 6142
rect 32732 6038 32788 6076
rect 32396 5908 32452 5918
rect 32396 5814 32452 5852
rect 32620 5684 32676 5694
rect 32620 5590 32676 5628
rect 32732 5682 32788 5694
rect 32732 5630 32734 5682
rect 32786 5630 32788 5682
rect 32732 5236 32788 5630
rect 32844 5572 32900 7422
rect 32956 6580 33012 6590
rect 32956 6486 33012 6524
rect 32844 5506 32900 5516
rect 32620 5012 32676 5022
rect 32620 4918 32676 4956
rect 32284 4274 32340 4284
rect 32172 3668 32228 3678
rect 32060 3666 32228 3668
rect 32060 3614 32174 3666
rect 32226 3614 32228 3666
rect 32060 3612 32228 3614
rect 32172 3602 32228 3612
rect 31836 3502 31838 3554
rect 31890 3502 31892 3554
rect 31836 3490 31892 3502
rect 32396 3556 32452 3566
rect 32732 3556 32788 5180
rect 32844 4564 32900 4574
rect 33068 4564 33124 7868
rect 33516 7812 33572 7822
rect 33516 5796 33572 7756
rect 33740 7698 33796 7980
rect 33740 7646 33742 7698
rect 33794 7646 33796 7698
rect 33740 7634 33796 7646
rect 33628 7476 33684 7486
rect 33628 7362 33684 7420
rect 33628 7310 33630 7362
rect 33682 7310 33684 7362
rect 33628 7298 33684 7310
rect 33964 7250 34020 7262
rect 33964 7198 33966 7250
rect 34018 7198 34020 7250
rect 33964 6692 34020 7198
rect 33964 6626 34020 6636
rect 33628 5796 33684 5806
rect 33516 5794 33684 5796
rect 33516 5742 33630 5794
rect 33682 5742 33684 5794
rect 33516 5740 33684 5742
rect 33628 5730 33684 5740
rect 32900 4508 33124 4564
rect 33180 5684 33236 5694
rect 32844 4226 32900 4508
rect 32844 4174 32846 4226
rect 32898 4174 32900 4226
rect 32844 4162 32900 4174
rect 33180 3666 33236 5628
rect 33740 5236 33796 5246
rect 33740 5142 33796 5180
rect 33180 3614 33182 3666
rect 33234 3614 33236 3666
rect 33180 3602 33236 3614
rect 33404 4564 33460 4574
rect 32396 3554 32788 3556
rect 32396 3502 32398 3554
rect 32450 3502 32788 3554
rect 32396 3500 32788 3502
rect 32396 3490 32452 3500
rect 32508 3332 32564 3342
rect 32508 3238 32564 3276
rect 31164 2482 31220 2492
rect 32060 1540 32116 1550
rect 32060 800 32116 1484
rect 33404 800 33460 4508
rect 33628 4228 33684 4238
rect 33628 4134 33684 4172
rect 34300 4116 34356 10108
rect 34524 9044 34580 10556
rect 34636 10498 34692 10510
rect 34636 10446 34638 10498
rect 34690 10446 34692 10498
rect 34636 10164 34692 10446
rect 34636 10098 34692 10108
rect 34636 9268 34692 9278
rect 34748 9268 34804 13580
rect 34972 13634 35028 13646
rect 34972 13582 34974 13634
rect 35026 13582 35028 13634
rect 34972 13412 35028 13582
rect 35420 13524 35476 14254
rect 35420 13458 35476 13468
rect 35532 13748 35588 13758
rect 34860 12180 34916 12190
rect 34860 11394 34916 12124
rect 34860 11342 34862 11394
rect 34914 11342 34916 11394
rect 34860 11172 34916 11342
rect 34972 11396 35028 13356
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13076 35252 13086
rect 35196 12982 35252 13020
rect 35532 12402 35588 13692
rect 35532 12350 35534 12402
rect 35586 12350 35588 12402
rect 35532 12338 35588 12350
rect 35084 12292 35140 12302
rect 35084 12198 35140 12236
rect 35308 12180 35364 12190
rect 35308 12086 35364 12124
rect 35532 11954 35588 11966
rect 35532 11902 35534 11954
rect 35586 11902 35588 11954
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11396 35140 11406
rect 34972 11394 35140 11396
rect 34972 11342 35086 11394
rect 35138 11342 35140 11394
rect 34972 11340 35140 11342
rect 35084 11330 35140 11340
rect 34860 11116 35028 11172
rect 34860 10948 34916 10958
rect 34860 10386 34916 10892
rect 34972 10836 35028 11116
rect 35532 10948 35588 11902
rect 35532 10882 35588 10892
rect 34972 10770 35028 10780
rect 35644 10724 35700 15148
rect 35756 13300 35812 16156
rect 35868 16100 35924 16604
rect 35980 16436 36036 17502
rect 35980 16370 36036 16380
rect 36092 17442 36148 17454
rect 36092 17390 36094 17442
rect 36146 17390 36148 17442
rect 35980 16100 36036 16110
rect 35868 16098 36036 16100
rect 35868 16046 35982 16098
rect 36034 16046 36036 16098
rect 35868 16044 36036 16046
rect 35980 16034 36036 16044
rect 36092 15876 36148 17390
rect 36204 17108 36260 18958
rect 36316 19012 36372 20132
rect 36428 19236 36484 22204
rect 36540 20468 36596 22540
rect 36652 21700 36708 23660
rect 36764 23042 36820 23054
rect 36764 22990 36766 23042
rect 36818 22990 36820 23042
rect 36764 22930 36820 22990
rect 37100 23044 37156 23054
rect 37100 22950 37156 22988
rect 36764 22878 36766 22930
rect 36818 22878 36820 22930
rect 36764 22866 36820 22878
rect 37436 22146 37492 22158
rect 37436 22094 37438 22146
rect 37490 22094 37492 22146
rect 37324 22036 37380 22046
rect 36652 21644 37044 21700
rect 36764 21474 36820 21486
rect 36764 21422 36766 21474
rect 36818 21422 36820 21474
rect 36652 20692 36708 20702
rect 36652 20598 36708 20636
rect 36540 20402 36596 20412
rect 36764 20188 36820 21422
rect 36988 20244 37044 21644
rect 37212 21474 37268 21486
rect 37212 21422 37214 21474
rect 37266 21422 37268 21474
rect 37212 21362 37268 21422
rect 37212 21310 37214 21362
rect 37266 21310 37268 21362
rect 37212 21298 37268 21310
rect 36764 20132 36932 20188
rect 36764 19906 36820 19918
rect 36764 19854 36766 19906
rect 36818 19854 36820 19906
rect 36764 19348 36820 19854
rect 36764 19282 36820 19292
rect 36428 19170 36484 19180
rect 36652 19012 36708 19022
rect 36316 19010 36820 19012
rect 36316 18958 36654 19010
rect 36706 18958 36820 19010
rect 36316 18956 36820 18958
rect 36652 18946 36708 18956
rect 36316 18450 36372 18462
rect 36316 18398 36318 18450
rect 36370 18398 36372 18450
rect 36316 18340 36372 18398
rect 36428 18340 36484 18350
rect 36316 18338 36484 18340
rect 36316 18286 36430 18338
rect 36482 18286 36484 18338
rect 36316 18284 36484 18286
rect 36428 18274 36484 18284
rect 36652 18340 36708 18350
rect 36540 18226 36596 18238
rect 36540 18174 36542 18226
rect 36594 18174 36596 18226
rect 36204 16772 36260 17052
rect 36316 17442 36372 17454
rect 36316 17390 36318 17442
rect 36370 17390 36372 17442
rect 36316 16996 36372 17390
rect 36540 17108 36596 18174
rect 36540 17042 36596 17052
rect 36652 18116 36708 18284
rect 36652 17442 36708 18060
rect 36652 17390 36654 17442
rect 36706 17390 36708 17442
rect 36316 16930 36372 16940
rect 36652 16884 36708 17390
rect 36652 16818 36708 16828
rect 36204 16716 36484 16772
rect 35868 15820 36148 15876
rect 36204 16436 36260 16446
rect 35868 15538 35924 15820
rect 36204 15764 36260 16380
rect 36316 16100 36372 16110
rect 36316 16006 36372 16044
rect 35868 15486 35870 15538
rect 35922 15486 35924 15538
rect 35868 15474 35924 15486
rect 36092 15708 36260 15764
rect 36316 15876 36372 15886
rect 36092 14418 36148 15708
rect 36316 15428 36372 15820
rect 36428 15538 36484 16716
rect 36540 16770 36596 16782
rect 36540 16718 36542 16770
rect 36594 16718 36596 16770
rect 36540 16212 36596 16718
rect 36764 16436 36820 18956
rect 36764 16370 36820 16380
rect 36876 18340 36932 20132
rect 36540 16146 36596 16156
rect 36540 15988 36596 15998
rect 36540 15894 36596 15932
rect 36652 15876 36708 15914
rect 36708 15820 36820 15876
rect 36652 15810 36708 15820
rect 36428 15486 36430 15538
rect 36482 15486 36484 15538
rect 36428 15474 36484 15486
rect 36652 15652 36708 15662
rect 36652 15538 36708 15596
rect 36652 15486 36654 15538
rect 36706 15486 36708 15538
rect 36652 15474 36708 15486
rect 36764 15540 36820 15820
rect 36764 15474 36820 15484
rect 36316 15296 36372 15372
rect 36428 15316 36484 15326
rect 36204 14642 36260 14654
rect 36204 14590 36206 14642
rect 36258 14590 36260 14642
rect 36204 14532 36260 14590
rect 36204 14466 36260 14476
rect 36092 14366 36094 14418
rect 36146 14366 36148 14418
rect 35980 13860 36036 13870
rect 35980 13766 36036 13804
rect 35868 13746 35924 13758
rect 35868 13694 35870 13746
rect 35922 13694 35924 13746
rect 35868 13524 35924 13694
rect 36092 13748 36148 14366
rect 36316 14306 36372 14318
rect 36316 14254 36318 14306
rect 36370 14254 36372 14306
rect 36204 13972 36260 13982
rect 36316 13972 36372 14254
rect 36204 13970 36372 13972
rect 36204 13918 36206 13970
rect 36258 13918 36372 13970
rect 36204 13916 36372 13918
rect 36204 13906 36260 13916
rect 36092 13692 36260 13748
rect 35868 13458 35924 13468
rect 35756 13244 35924 13300
rect 35756 13076 35812 13086
rect 35756 12962 35812 13020
rect 35756 12910 35758 12962
rect 35810 12910 35812 12962
rect 35756 12898 35812 12910
rect 35868 12850 35924 13244
rect 35868 12798 35870 12850
rect 35922 12798 35924 12850
rect 35868 12292 35924 12798
rect 36092 12852 36148 12862
rect 36092 12758 36148 12796
rect 36204 12628 36260 13692
rect 36204 12562 36260 12572
rect 36316 13300 36372 13310
rect 35868 12226 35924 12236
rect 35756 12178 35812 12190
rect 35756 12126 35758 12178
rect 35810 12126 35812 12178
rect 35756 12068 35812 12126
rect 35756 12002 35812 12012
rect 36092 12178 36148 12190
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 36092 11844 36148 12126
rect 36316 11844 36372 13244
rect 36428 12740 36484 15260
rect 36540 14306 36596 14318
rect 36540 14254 36542 14306
rect 36594 14254 36596 14306
rect 36540 13972 36596 14254
rect 36652 13972 36708 13982
rect 36540 13970 36708 13972
rect 36540 13918 36654 13970
rect 36706 13918 36708 13970
rect 36540 13916 36708 13918
rect 36652 13906 36708 13916
rect 36540 13748 36596 13758
rect 36540 12852 36596 13692
rect 36652 13524 36708 13534
rect 36652 13186 36708 13468
rect 36652 13134 36654 13186
rect 36706 13134 36708 13186
rect 36652 13122 36708 13134
rect 36652 12852 36708 12862
rect 36540 12850 36708 12852
rect 36540 12798 36654 12850
rect 36706 12798 36708 12850
rect 36540 12796 36708 12798
rect 36652 12786 36708 12796
rect 36764 12852 36820 12862
rect 36764 12758 36820 12796
rect 36428 12684 36596 12740
rect 36428 12516 36484 12526
rect 36428 12402 36484 12460
rect 36428 12350 36430 12402
rect 36482 12350 36484 12402
rect 36428 12338 36484 12350
rect 36092 11788 36372 11844
rect 36540 11788 36596 12684
rect 36652 12404 36708 12414
rect 36652 12310 36708 12348
rect 36764 12292 36820 12302
rect 36764 12198 36820 12236
rect 36092 11620 36148 11630
rect 36092 11394 36148 11564
rect 36092 11342 36094 11394
rect 36146 11342 36148 11394
rect 36092 11330 36148 11342
rect 36092 11170 36148 11182
rect 36092 11118 36094 11170
rect 36146 11118 36148 11170
rect 36092 11060 36148 11118
rect 36092 10994 36148 11004
rect 36316 10948 36372 11788
rect 36316 10882 36372 10892
rect 36428 11732 36596 11788
rect 35980 10836 36036 10846
rect 35980 10742 36036 10780
rect 35868 10724 35924 10734
rect 35644 10722 35924 10724
rect 35644 10670 35870 10722
rect 35922 10670 35924 10722
rect 35644 10668 35924 10670
rect 34972 10612 35028 10622
rect 34972 10518 35028 10556
rect 35308 10612 35364 10622
rect 34860 10334 34862 10386
rect 34914 10334 34916 10386
rect 34860 10164 34916 10334
rect 35308 10388 35364 10556
rect 35420 10612 35476 10622
rect 35420 10610 35588 10612
rect 35420 10558 35422 10610
rect 35474 10558 35588 10610
rect 35420 10556 35588 10558
rect 35420 10546 35476 10556
rect 35308 10322 35364 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 34860 10108 35140 10164
rect 35196 10154 35460 10164
rect 34636 9266 34804 9268
rect 34636 9214 34638 9266
rect 34690 9214 34804 9266
rect 34636 9212 34804 9214
rect 34636 9202 34692 9212
rect 34748 9044 34804 9054
rect 34524 8988 34692 9044
rect 34524 7474 34580 7486
rect 34524 7422 34526 7474
rect 34578 7422 34580 7474
rect 34524 5124 34580 7422
rect 34636 7476 34692 8988
rect 34748 8950 34804 8988
rect 34860 8932 34916 8942
rect 34860 8838 34916 8876
rect 34972 8820 35028 8830
rect 34860 7476 34916 7486
rect 34636 7420 34860 7476
rect 34860 7382 34916 7420
rect 34972 6804 35028 8764
rect 35084 7252 35140 10108
rect 35308 9940 35364 9950
rect 35308 9846 35364 9884
rect 35532 9380 35588 10556
rect 35868 10052 35924 10668
rect 35980 10612 36036 10622
rect 35980 10386 36036 10556
rect 35980 10334 35982 10386
rect 36034 10334 36036 10386
rect 35980 10164 36036 10334
rect 35980 10098 36036 10108
rect 36092 10388 36148 10398
rect 35868 9986 35924 9996
rect 36092 9940 36148 10332
rect 36428 10388 36484 11732
rect 36764 11508 36820 11518
rect 36764 11284 36820 11452
rect 36764 11218 36820 11228
rect 36652 11172 36708 11182
rect 36428 10322 36484 10332
rect 36540 10724 36596 10734
rect 36540 10498 36596 10668
rect 36540 10446 36542 10498
rect 36594 10446 36596 10498
rect 36540 10276 36596 10446
rect 36540 10210 36596 10220
rect 36652 10050 36708 11116
rect 36652 9998 36654 10050
rect 36706 9998 36708 10050
rect 36652 9986 36708 9998
rect 36764 10388 36820 10398
rect 35980 9884 36148 9940
rect 36764 9938 36820 10332
rect 36764 9886 36766 9938
rect 36818 9886 36820 9938
rect 35980 9714 36036 9884
rect 36764 9874 36820 9886
rect 36204 9828 36260 9838
rect 35980 9662 35982 9714
rect 36034 9662 36036 9714
rect 35756 9604 35812 9614
rect 35532 9314 35588 9324
rect 35644 9602 35812 9604
rect 35644 9550 35758 9602
rect 35810 9550 35812 9602
rect 35644 9548 35812 9550
rect 35420 9042 35476 9054
rect 35420 8990 35422 9042
rect 35474 8990 35476 9042
rect 35420 8820 35476 8990
rect 35532 8932 35588 8942
rect 35532 8838 35588 8876
rect 35420 8754 35476 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35532 8370 35588 8382
rect 35532 8318 35534 8370
rect 35586 8318 35588 8370
rect 35532 7924 35588 8318
rect 35644 8260 35700 9548
rect 35756 9538 35812 9548
rect 35980 9492 36036 9662
rect 36092 9716 36148 9726
rect 36204 9716 36260 9772
rect 36092 9714 36260 9716
rect 36092 9662 36094 9714
rect 36146 9662 36260 9714
rect 36092 9660 36260 9662
rect 36092 9650 36148 9660
rect 35980 9426 36036 9436
rect 36652 9156 36708 9166
rect 36540 9100 36652 9156
rect 36316 8930 36372 8942
rect 36316 8878 36318 8930
rect 36370 8878 36372 8930
rect 35644 8194 35700 8204
rect 35756 8818 35812 8830
rect 35756 8766 35758 8818
rect 35810 8766 35812 8818
rect 35756 8036 35812 8766
rect 36092 8260 36148 8270
rect 35756 7970 35812 7980
rect 35980 8258 36148 8260
rect 35980 8206 36094 8258
rect 36146 8206 36148 8258
rect 35980 8204 36148 8206
rect 35532 7858 35588 7868
rect 35420 7812 35476 7822
rect 35420 7588 35476 7756
rect 35644 7700 35700 7710
rect 35980 7700 36036 8204
rect 36092 8194 36148 8204
rect 36316 8260 36372 8878
rect 36428 8372 36484 8382
rect 36428 8278 36484 8316
rect 36316 8194 36372 8204
rect 36540 8258 36596 9100
rect 36652 9062 36708 9100
rect 36876 8932 36932 18284
rect 36988 15148 37044 20188
rect 37212 20020 37268 20030
rect 37100 19908 37156 19918
rect 37100 19814 37156 19852
rect 37100 18340 37156 18350
rect 37100 18246 37156 18284
rect 37212 18226 37268 19964
rect 37324 19794 37380 21980
rect 37436 21924 37492 22094
rect 37436 21858 37492 21868
rect 37548 21810 37604 23996
rect 37772 23716 37828 23726
rect 38220 23716 38276 23726
rect 37772 23714 38276 23716
rect 37772 23662 37774 23714
rect 37826 23662 38222 23714
rect 38274 23662 38276 23714
rect 37772 23660 38276 23662
rect 37772 23650 37828 23660
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 37884 22372 37940 22382
rect 37884 22036 37940 22316
rect 37884 21970 37940 21980
rect 37548 21758 37550 21810
rect 37602 21758 37604 21810
rect 37436 20804 37492 20814
rect 37436 20710 37492 20748
rect 37548 20188 37604 21758
rect 37996 21474 38052 21486
rect 37996 21422 37998 21474
rect 38050 21422 38052 21474
rect 37996 20916 38052 21422
rect 37996 20850 38052 20860
rect 38108 21362 38164 21374
rect 38108 21310 38110 21362
rect 38162 21310 38164 21362
rect 37884 20578 37940 20590
rect 37884 20526 37886 20578
rect 37938 20526 37940 20578
rect 37548 20132 37828 20188
rect 37324 19742 37326 19794
rect 37378 19742 37380 19794
rect 37324 19730 37380 19742
rect 37548 19906 37604 19918
rect 37548 19854 37550 19906
rect 37602 19854 37604 19906
rect 37548 19684 37604 19854
rect 37548 19618 37604 19628
rect 37436 19458 37492 19470
rect 37436 19406 37438 19458
rect 37490 19406 37492 19458
rect 37436 19010 37492 19406
rect 37436 18958 37438 19010
rect 37490 18958 37492 19010
rect 37436 18900 37492 18958
rect 37436 18834 37492 18844
rect 37548 19236 37604 19246
rect 37212 18174 37214 18226
rect 37266 18174 37268 18226
rect 37212 18004 37268 18174
rect 37212 17938 37268 17948
rect 37548 17780 37604 19180
rect 37772 18452 37828 20132
rect 37884 20020 37940 20526
rect 37884 19954 37940 19964
rect 37996 20244 38052 20254
rect 37996 20018 38052 20188
rect 37996 19966 37998 20018
rect 38050 19966 38052 20018
rect 37996 19954 38052 19966
rect 37884 19794 37940 19806
rect 37884 19742 37886 19794
rect 37938 19742 37940 19794
rect 37884 19346 37940 19742
rect 37884 19294 37886 19346
rect 37938 19294 37940 19346
rect 37884 19282 37940 19294
rect 37996 19796 38052 19806
rect 37772 18386 37828 18396
rect 37660 18340 37716 18350
rect 37660 18246 37716 18284
rect 37884 18228 37940 18238
rect 37996 18228 38052 19740
rect 38108 19236 38164 21310
rect 38108 19170 38164 19180
rect 37884 18226 38052 18228
rect 37884 18174 37886 18226
rect 37938 18174 38052 18226
rect 37884 18172 38052 18174
rect 38108 19012 38164 19022
rect 38220 19012 38276 23660
rect 38332 23042 38388 23054
rect 38332 22990 38334 23042
rect 38386 22990 38388 23042
rect 38332 22484 38388 22990
rect 38332 22418 38388 22428
rect 38444 22484 38500 24780
rect 41580 24610 41636 24622
rect 41580 24558 41582 24610
rect 41634 24558 41636 24610
rect 39452 23828 39508 23838
rect 39452 23734 39508 23772
rect 38668 23714 38724 23726
rect 38668 23662 38670 23714
rect 38722 23662 38724 23714
rect 38556 22484 38612 22494
rect 38444 22482 38612 22484
rect 38444 22430 38558 22482
rect 38610 22430 38612 22482
rect 38444 22428 38612 22430
rect 38332 22260 38388 22270
rect 38444 22260 38500 22428
rect 38556 22418 38612 22428
rect 38668 22484 38724 23662
rect 39116 23714 39172 23726
rect 39116 23662 39118 23714
rect 39170 23662 39172 23714
rect 38668 22418 38724 22428
rect 38780 23042 38836 23054
rect 38780 22990 38782 23042
rect 38834 22990 38836 23042
rect 38780 22372 38836 22990
rect 39004 22708 39060 22718
rect 38780 22306 38836 22316
rect 38892 22482 38948 22494
rect 38892 22430 38894 22482
rect 38946 22430 38948 22482
rect 38892 22370 38948 22430
rect 38892 22318 38894 22370
rect 38946 22318 38948 22370
rect 38892 22306 38948 22318
rect 38332 22258 38500 22260
rect 38332 22206 38334 22258
rect 38386 22206 38500 22258
rect 38332 22204 38500 22206
rect 38332 22194 38388 22204
rect 38892 22148 38948 22158
rect 38892 21810 38948 22092
rect 38892 21758 38894 21810
rect 38946 21758 38948 21810
rect 38892 21746 38948 21758
rect 38332 21700 38388 21710
rect 38332 20578 38388 21644
rect 38444 21474 38500 21486
rect 38444 21422 38446 21474
rect 38498 21422 38500 21474
rect 38444 21364 38500 21422
rect 38444 21298 38500 21308
rect 38780 21028 38836 21038
rect 38780 20914 38836 20972
rect 38780 20862 38782 20914
rect 38834 20862 38836 20914
rect 38780 20850 38836 20862
rect 38332 20526 38334 20578
rect 38386 20526 38388 20578
rect 38332 19458 38388 20526
rect 38444 19908 38500 19918
rect 38444 19814 38500 19852
rect 38892 19906 38948 19918
rect 38892 19854 38894 19906
rect 38946 19854 38948 19906
rect 38332 19406 38334 19458
rect 38386 19406 38388 19458
rect 38332 19394 38388 19406
rect 38164 18956 38276 19012
rect 38332 19010 38388 19022
rect 38332 18958 38334 19010
rect 38386 18958 38388 19010
rect 38108 18338 38164 18956
rect 38108 18286 38110 18338
rect 38162 18286 38164 18338
rect 37548 17724 37828 17780
rect 37548 17556 37604 17566
rect 37436 17554 37604 17556
rect 37436 17502 37550 17554
rect 37602 17502 37604 17554
rect 37436 17500 37604 17502
rect 37100 17108 37156 17118
rect 37100 17014 37156 17052
rect 37324 17108 37380 17118
rect 37324 17014 37380 17052
rect 37324 16884 37380 16894
rect 37212 16770 37268 16782
rect 37212 16718 37214 16770
rect 37266 16718 37268 16770
rect 37212 15988 37268 16718
rect 37212 15922 37268 15932
rect 37212 15764 37268 15774
rect 37212 15538 37268 15708
rect 37212 15486 37214 15538
rect 37266 15486 37268 15538
rect 37212 15474 37268 15486
rect 37100 15428 37156 15438
rect 37100 15334 37156 15372
rect 36988 15092 37268 15148
rect 37100 14644 37156 14654
rect 36988 13524 37044 13534
rect 36988 13430 37044 13468
rect 37100 11508 37156 14588
rect 37212 14420 37268 15092
rect 37324 14644 37380 16828
rect 37436 16212 37492 17500
rect 37548 17490 37604 17500
rect 37660 17442 37716 17454
rect 37660 17390 37662 17442
rect 37714 17390 37716 17442
rect 37660 16882 37716 17390
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 37660 16818 37716 16830
rect 37772 16436 37828 17724
rect 37436 16098 37492 16156
rect 37436 16046 37438 16098
rect 37490 16046 37492 16098
rect 37436 15652 37492 16046
rect 37436 15586 37492 15596
rect 37548 16380 37828 16436
rect 37436 15428 37492 15438
rect 37436 15334 37492 15372
rect 37548 15148 37604 16380
rect 37660 16210 37716 16222
rect 37660 16158 37662 16210
rect 37714 16158 37716 16210
rect 37660 16100 37716 16158
rect 37660 16034 37716 16044
rect 37772 15874 37828 15886
rect 37772 15822 37774 15874
rect 37826 15822 37828 15874
rect 37772 15764 37828 15822
rect 37772 15698 37828 15708
rect 37884 15540 37940 18172
rect 38108 17668 38164 18286
rect 38108 17602 38164 17612
rect 38108 17444 38164 17454
rect 38108 17350 38164 17388
rect 38220 17442 38276 17454
rect 38220 17390 38222 17442
rect 38274 17390 38276 17442
rect 38220 17220 38276 17390
rect 37996 17164 38276 17220
rect 38332 17220 38388 18958
rect 38780 19010 38836 19022
rect 38780 18958 38782 19010
rect 38834 18958 38836 19010
rect 38780 18900 38836 18958
rect 38780 18834 38836 18844
rect 38556 18338 38612 18350
rect 38556 18286 38558 18338
rect 38610 18286 38612 18338
rect 38556 18226 38612 18286
rect 38556 18174 38558 18226
rect 38610 18174 38612 18226
rect 38556 18162 38612 18174
rect 38892 18116 38948 19854
rect 39004 18450 39060 22652
rect 39116 19908 39172 23662
rect 40236 23716 40292 23726
rect 40236 23622 40292 23660
rect 40684 23714 40740 23726
rect 40684 23662 40686 23714
rect 40738 23662 40740 23714
rect 40684 23604 40740 23662
rect 40684 23538 40740 23548
rect 41356 23714 41412 23726
rect 41356 23662 41358 23714
rect 41410 23662 41412 23714
rect 41244 23492 41300 23502
rect 39676 23268 39732 23278
rect 39676 23174 39732 23212
rect 39228 23044 39284 23054
rect 39228 22950 39284 22988
rect 40236 23042 40292 23054
rect 40236 22990 40238 23042
rect 40290 22990 40292 23042
rect 39900 22596 39956 22606
rect 39676 22036 39732 22046
rect 39340 21812 39396 21822
rect 39340 21476 39396 21756
rect 39340 21382 39396 21420
rect 39228 20580 39284 20590
rect 39228 20486 39284 20524
rect 39340 20132 39396 20142
rect 39340 20038 39396 20076
rect 39116 19842 39172 19852
rect 39676 19458 39732 21980
rect 39900 21924 39956 22540
rect 40012 22258 40068 22270
rect 40012 22206 40014 22258
rect 40066 22206 40068 22258
rect 40012 22036 40068 22206
rect 40012 21970 40068 21980
rect 39900 21476 39956 21868
rect 40236 21700 40292 22990
rect 40684 23042 40740 23054
rect 40684 22990 40686 23042
rect 40738 22990 40740 23042
rect 40572 22148 40628 22158
rect 40572 22054 40628 22092
rect 40236 21634 40292 21644
rect 40460 21812 40516 21822
rect 40012 21476 40068 21486
rect 40460 21476 40516 21756
rect 39900 21474 40068 21476
rect 39900 21422 40014 21474
rect 40066 21422 40068 21474
rect 39900 21420 40068 21422
rect 39788 19906 39844 19918
rect 39788 19854 39790 19906
rect 39842 19854 39844 19906
rect 39788 19572 39844 19854
rect 39788 19506 39844 19516
rect 39676 19406 39678 19458
rect 39730 19406 39732 19458
rect 39676 19394 39732 19406
rect 39676 19124 39732 19134
rect 39676 19030 39732 19068
rect 39228 19012 39284 19022
rect 39228 18918 39284 18956
rect 39900 18900 39956 21420
rect 40012 21410 40068 21420
rect 40348 21474 40516 21476
rect 40348 21422 40462 21474
rect 40514 21422 40516 21474
rect 40348 21420 40516 21422
rect 40348 20692 40404 21420
rect 40460 21410 40516 21420
rect 40124 20636 40404 20692
rect 40012 20578 40068 20590
rect 40012 20526 40014 20578
rect 40066 20526 40068 20578
rect 40012 20468 40068 20526
rect 40012 20402 40068 20412
rect 39900 18834 39956 18844
rect 40012 19012 40068 19022
rect 39004 18398 39006 18450
rect 39058 18398 39060 18450
rect 39004 18386 39060 18398
rect 39452 18452 39508 18462
rect 39452 18358 39508 18396
rect 39900 18338 39956 18350
rect 39900 18286 39902 18338
rect 39954 18286 39956 18338
rect 39900 18228 39956 18286
rect 39900 18162 39956 18172
rect 38892 18050 38948 18060
rect 38780 17666 38836 17678
rect 38780 17614 38782 17666
rect 38834 17614 38836 17666
rect 38444 17444 38500 17454
rect 38444 17350 38500 17388
rect 38332 17164 38500 17220
rect 37996 16884 38052 17164
rect 38332 16996 38388 17006
rect 38332 16902 38388 16940
rect 37996 15986 38052 16828
rect 37996 15934 37998 15986
rect 38050 15934 38052 15986
rect 37996 15922 38052 15934
rect 37324 14578 37380 14588
rect 37436 15092 37604 15148
rect 37660 15484 37940 15540
rect 37212 14364 37380 14420
rect 37212 13860 37268 13870
rect 37212 13766 37268 13804
rect 37324 13300 37380 14364
rect 37436 14308 37492 15092
rect 37660 14418 37716 15484
rect 38332 15428 38388 15438
rect 38332 15334 38388 15372
rect 37660 14366 37662 14418
rect 37714 14366 37716 14418
rect 37436 14242 37492 14252
rect 37548 14306 37604 14318
rect 37548 14254 37550 14306
rect 37602 14254 37604 14306
rect 37324 13234 37380 13244
rect 37548 13972 37604 14254
rect 37324 12852 37380 12862
rect 37100 11442 37156 11452
rect 37212 12516 37268 12526
rect 37100 10500 37156 10510
rect 37100 10406 37156 10444
rect 37100 10276 37156 10286
rect 36876 8866 36932 8876
rect 36988 9492 37044 9502
rect 36540 8206 36542 8258
rect 36594 8206 36596 8258
rect 36540 8194 36596 8206
rect 36764 8148 36820 8158
rect 36764 8146 36932 8148
rect 36764 8094 36766 8146
rect 36818 8094 36932 8146
rect 36764 8092 36932 8094
rect 36764 8082 36820 8092
rect 36316 8036 36372 8046
rect 36316 7942 36372 7980
rect 35644 7698 36036 7700
rect 35644 7646 35646 7698
rect 35698 7646 36036 7698
rect 35644 7644 36036 7646
rect 36092 7924 36148 7934
rect 35644 7634 35700 7644
rect 35532 7588 35588 7598
rect 35420 7586 35588 7588
rect 35420 7534 35534 7586
rect 35586 7534 35588 7586
rect 35420 7532 35588 7534
rect 35532 7522 35588 7532
rect 36092 7586 36148 7868
rect 36764 7812 36820 7822
rect 36092 7534 36094 7586
rect 36146 7534 36148 7586
rect 36092 7522 36148 7534
rect 36652 7698 36708 7710
rect 36652 7646 36654 7698
rect 36706 7646 36708 7698
rect 35308 7364 35364 7374
rect 35308 7270 35364 7308
rect 36316 7364 36372 7374
rect 36316 7270 36372 7308
rect 35084 7158 35140 7196
rect 36540 7252 36596 7262
rect 36540 7158 36596 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6804 35140 6814
rect 34972 6802 35140 6804
rect 34972 6750 35086 6802
rect 35138 6750 35140 6802
rect 34972 6748 35140 6750
rect 35084 6020 35140 6748
rect 36652 6690 36708 7646
rect 36764 7476 36820 7756
rect 36764 7382 36820 7420
rect 36652 6638 36654 6690
rect 36706 6638 36708 6690
rect 36652 6626 36708 6638
rect 35084 5954 35140 5964
rect 35980 6578 36036 6590
rect 35980 6526 35982 6578
rect 36034 6526 36036 6578
rect 35980 6468 36036 6526
rect 35980 6020 36036 6412
rect 36204 6466 36260 6478
rect 36204 6414 36206 6466
rect 36258 6414 36260 6466
rect 36204 6356 36260 6414
rect 36204 6290 36260 6300
rect 36316 6466 36372 6478
rect 36316 6414 36318 6466
rect 36370 6414 36372 6466
rect 35980 5954 36036 5964
rect 35756 5796 35812 5806
rect 36316 5796 36372 6414
rect 36428 6466 36484 6478
rect 36428 6414 36430 6466
rect 36482 6414 36484 6466
rect 36428 6132 36484 6414
rect 36428 6076 36596 6132
rect 35756 5702 35812 5740
rect 35980 5740 36372 5796
rect 36428 5906 36484 5918
rect 36428 5854 36430 5906
rect 36482 5854 36484 5906
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35756 5460 35812 5470
rect 35756 5346 35812 5404
rect 35756 5294 35758 5346
rect 35810 5294 35812 5346
rect 35756 5282 35812 5294
rect 35868 5348 35924 5358
rect 35868 5254 35924 5292
rect 34524 5058 34580 5068
rect 34972 5010 35028 5022
rect 34972 4958 34974 5010
rect 35026 4958 35028 5010
rect 34972 4564 35028 4958
rect 34972 4498 35028 4508
rect 35756 4452 35812 4462
rect 35980 4452 36036 5740
rect 36204 5572 36260 5582
rect 36092 5124 36148 5134
rect 36092 5030 36148 5068
rect 36204 4898 36260 5516
rect 36316 5124 36372 5134
rect 36316 5030 36372 5068
rect 36204 4846 36206 4898
rect 36258 4846 36260 4898
rect 36204 4834 36260 4846
rect 35756 4450 36036 4452
rect 35756 4398 35758 4450
rect 35810 4398 36036 4450
rect 35756 4396 36036 4398
rect 35756 4386 35812 4396
rect 36428 4340 36484 5854
rect 36428 4246 36484 4284
rect 34300 4050 34356 4060
rect 35532 4116 35588 4126
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35532 3778 35588 4060
rect 35532 3726 35534 3778
rect 35586 3726 35588 3778
rect 35532 3714 35588 3726
rect 35756 3780 35812 3790
rect 35756 3686 35812 3724
rect 35868 3668 35924 3678
rect 35868 3574 35924 3612
rect 35308 3554 35364 3566
rect 35308 3502 35310 3554
rect 35362 3502 35364 3554
rect 34524 3442 34580 3454
rect 34524 3390 34526 3442
rect 34578 3390 34580 3442
rect 34524 1540 34580 3390
rect 34524 1474 34580 1484
rect 34748 3444 34804 3454
rect 34748 2436 34804 3388
rect 35308 2660 35364 3502
rect 35420 3330 35476 3342
rect 35420 3278 35422 3330
rect 35474 3278 35476 3330
rect 35420 3220 35476 3278
rect 35420 2884 35476 3164
rect 36540 3108 36596 6076
rect 36876 6020 36932 8092
rect 36988 7812 37044 9436
rect 36988 7746 37044 7756
rect 36876 5954 36932 5964
rect 36988 7474 37044 7486
rect 36988 7422 36990 7474
rect 37042 7422 37044 7474
rect 36988 5124 37044 7422
rect 37100 7364 37156 10220
rect 37212 7588 37268 12460
rect 37324 12290 37380 12796
rect 37548 12516 37604 13916
rect 37660 13076 37716 14366
rect 37772 15202 37828 15214
rect 37772 15150 37774 15202
rect 37826 15150 37828 15202
rect 37772 14084 37828 15150
rect 38108 14308 38164 14318
rect 38108 14214 38164 14252
rect 38444 14196 38500 17164
rect 38668 17108 38724 17118
rect 38668 17014 38724 17052
rect 38556 16882 38612 16894
rect 38556 16830 38558 16882
rect 38610 16830 38612 16882
rect 38556 15874 38612 16830
rect 38556 15822 38558 15874
rect 38610 15822 38612 15874
rect 38556 15428 38612 15822
rect 38556 15362 38612 15372
rect 38668 16436 38724 16446
rect 38668 15314 38724 16380
rect 38780 16210 38836 17614
rect 39228 17554 39284 17566
rect 39228 17502 39230 17554
rect 39282 17502 39284 17554
rect 39004 17444 39060 17454
rect 39004 16884 39060 17388
rect 38780 16158 38782 16210
rect 38834 16158 38836 16210
rect 38780 16146 38836 16158
rect 38892 16882 39060 16884
rect 38892 16830 39006 16882
rect 39058 16830 39060 16882
rect 38892 16828 39060 16830
rect 38780 15988 38836 15998
rect 38892 15988 38948 16828
rect 39004 16818 39060 16828
rect 39116 16100 39172 16110
rect 39116 16006 39172 16044
rect 38780 15986 38892 15988
rect 38780 15934 38782 15986
rect 38834 15934 38892 15986
rect 38780 15932 38892 15934
rect 38780 15922 38836 15932
rect 38892 15856 38948 15932
rect 38668 15262 38670 15314
rect 38722 15262 38724 15314
rect 38668 15148 38724 15262
rect 38780 15316 38836 15326
rect 38780 15222 38836 15260
rect 38892 15316 38948 15326
rect 39228 15316 39284 17502
rect 39340 17444 39396 17454
rect 39340 17350 39396 17388
rect 40012 17442 40068 18956
rect 40124 18788 40180 20636
rect 40460 20578 40516 20590
rect 40460 20526 40462 20578
rect 40514 20526 40516 20578
rect 40348 19908 40404 19918
rect 40236 19458 40292 19470
rect 40236 19406 40238 19458
rect 40290 19406 40292 19458
rect 40236 19346 40292 19406
rect 40236 19294 40238 19346
rect 40290 19294 40292 19346
rect 40236 18900 40292 19294
rect 40348 19012 40404 19852
rect 40460 19796 40516 20526
rect 40460 19730 40516 19740
rect 40684 19348 40740 22990
rect 41020 22146 41076 22158
rect 41020 22094 41022 22146
rect 41074 22094 41076 22146
rect 41020 21924 41076 22094
rect 41020 21858 41076 21868
rect 41244 20914 41300 23436
rect 41356 22596 41412 23662
rect 41580 23156 41636 24558
rect 43148 24500 43204 24510
rect 42476 24164 42532 24174
rect 41580 23090 41636 23100
rect 41804 23714 41860 23726
rect 41804 23662 41806 23714
rect 41858 23662 41860 23714
rect 41468 23044 41524 23054
rect 41468 22950 41524 22988
rect 41356 22530 41412 22540
rect 41692 22146 41748 22158
rect 41692 22094 41694 22146
rect 41746 22094 41748 22146
rect 41692 21924 41748 22094
rect 41692 21858 41748 21868
rect 41804 21812 41860 23662
rect 42028 23268 42084 23278
rect 42028 23174 42084 23212
rect 42364 23268 42420 23278
rect 42140 22484 42196 22494
rect 42028 22146 42084 22158
rect 42028 22094 42030 22146
rect 42082 22094 42084 22146
rect 42028 22036 42084 22094
rect 41804 21746 41860 21756
rect 41916 21980 42084 22036
rect 41468 21476 41524 21486
rect 41244 20862 41246 20914
rect 41298 20862 41300 20914
rect 40684 19282 40740 19292
rect 40796 19906 40852 19918
rect 40796 19854 40798 19906
rect 40850 19854 40852 19906
rect 40684 19012 40740 19022
rect 40796 19012 40852 19854
rect 41244 19458 41300 20862
rect 41244 19406 41246 19458
rect 41298 19406 41300 19458
rect 41244 19394 41300 19406
rect 41356 21474 41524 21476
rect 41356 21422 41470 21474
rect 41522 21422 41524 21474
rect 41356 21420 41524 21422
rect 41356 19460 41412 21420
rect 41468 21410 41524 21420
rect 41916 21476 41972 21980
rect 42028 21812 42084 21822
rect 42140 21812 42196 22428
rect 42028 21810 42196 21812
rect 42028 21758 42030 21810
rect 42082 21758 42196 21810
rect 42028 21756 42196 21758
rect 42028 21746 42084 21756
rect 41580 20916 41636 20926
rect 41468 19908 41524 19918
rect 41468 19814 41524 19852
rect 41356 19394 41412 19404
rect 41356 19236 41412 19246
rect 41244 19012 41300 19022
rect 40348 18956 40516 19012
rect 40236 18844 40404 18900
rect 40124 18732 40292 18788
rect 40012 17390 40014 17442
rect 40066 17390 40068 17442
rect 40012 17220 40068 17390
rect 40012 17154 40068 17164
rect 40124 17780 40180 17790
rect 39564 16994 39620 17006
rect 39564 16942 39566 16994
rect 39618 16942 39620 16994
rect 39340 16884 39396 16894
rect 39340 16790 39396 16828
rect 39564 16436 39620 16942
rect 39788 16996 39844 17006
rect 39676 16884 39732 16894
rect 39676 16790 39732 16828
rect 39564 16380 39732 16436
rect 39564 16212 39620 16222
rect 39564 16118 39620 16156
rect 38892 15314 39284 15316
rect 38892 15262 38894 15314
rect 38946 15262 39284 15314
rect 38892 15260 39284 15262
rect 39340 16100 39396 16110
rect 38668 15092 38836 15148
rect 38780 14530 38836 15092
rect 38892 14868 38948 15260
rect 39340 15148 39396 16044
rect 39452 15988 39508 15998
rect 39452 15426 39508 15932
rect 39676 15540 39732 16380
rect 39788 15986 39844 16940
rect 39900 16436 39956 16446
rect 39900 16322 39956 16380
rect 39900 16270 39902 16322
rect 39954 16270 39956 16322
rect 39900 16258 39956 16270
rect 39788 15934 39790 15986
rect 39842 15934 39844 15986
rect 39788 15922 39844 15934
rect 39900 15876 39956 15886
rect 39788 15540 39844 15550
rect 39676 15538 39844 15540
rect 39676 15486 39790 15538
rect 39842 15486 39844 15538
rect 39676 15484 39844 15486
rect 39788 15474 39844 15484
rect 39452 15374 39454 15426
rect 39506 15374 39508 15426
rect 39452 15362 39508 15374
rect 39564 15428 39620 15438
rect 39564 15148 39620 15372
rect 38892 14802 38948 14812
rect 39004 15092 39396 15148
rect 39452 15092 39620 15148
rect 38780 14478 38782 14530
rect 38834 14478 38836 14530
rect 38780 14466 38836 14478
rect 38444 14130 38500 14140
rect 38892 14306 38948 14318
rect 38892 14254 38894 14306
rect 38946 14254 38948 14306
rect 37772 14018 37828 14028
rect 37660 13010 37716 13020
rect 37772 13860 37828 13870
rect 37772 13074 37828 13804
rect 38332 13860 38388 13870
rect 38332 13766 38388 13804
rect 38220 13748 38276 13758
rect 38108 13524 38164 13534
rect 38108 13430 38164 13468
rect 37772 13022 37774 13074
rect 37826 13022 37828 13074
rect 37772 13010 37828 13022
rect 38220 12962 38276 13692
rect 38892 13746 38948 14254
rect 38892 13694 38894 13746
rect 38946 13694 38948 13746
rect 38444 13636 38500 13646
rect 38892 13636 38948 13694
rect 38444 13634 38948 13636
rect 38444 13582 38446 13634
rect 38498 13582 38948 13634
rect 38444 13580 38948 13582
rect 38444 13570 38500 13580
rect 39004 13076 39060 15092
rect 39116 14420 39172 14430
rect 39116 14326 39172 14364
rect 39452 13970 39508 15092
rect 39900 14644 39956 15820
rect 39900 14578 39956 14588
rect 40012 15764 40068 15774
rect 39564 14420 39620 14430
rect 39564 14326 39620 14364
rect 39900 14420 39956 14430
rect 39900 14326 39956 14364
rect 39452 13918 39454 13970
rect 39506 13918 39508 13970
rect 39452 13906 39508 13918
rect 39564 13972 39620 13982
rect 39564 13878 39620 13916
rect 40012 13970 40068 15708
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 40012 13906 40068 13918
rect 39676 13860 39732 13870
rect 39340 13748 39396 13758
rect 39340 13746 39508 13748
rect 39340 13694 39342 13746
rect 39394 13694 39508 13746
rect 39340 13692 39508 13694
rect 39340 13682 39396 13692
rect 39340 13412 39396 13422
rect 38892 13020 39060 13076
rect 39116 13076 39172 13086
rect 38556 12964 38612 12974
rect 38220 12910 38222 12962
rect 38274 12910 38276 12962
rect 38220 12898 38276 12910
rect 38332 12908 38556 12964
rect 37660 12852 37716 12862
rect 37996 12852 38052 12862
rect 37660 12758 37716 12796
rect 37772 12850 38052 12852
rect 37772 12798 37998 12850
rect 38050 12798 38052 12850
rect 37772 12796 38052 12798
rect 37772 12740 37828 12796
rect 37996 12786 38052 12796
rect 38108 12852 38164 12862
rect 37772 12674 37828 12684
rect 37548 12460 37940 12516
rect 37436 12404 37492 12414
rect 37436 12402 37604 12404
rect 37436 12350 37438 12402
rect 37490 12350 37604 12402
rect 37436 12348 37604 12350
rect 37436 12338 37492 12348
rect 37324 12238 37326 12290
rect 37378 12238 37380 12290
rect 37324 12226 37380 12238
rect 37436 11954 37492 11966
rect 37436 11902 37438 11954
rect 37490 11902 37492 11954
rect 37436 11844 37492 11902
rect 37436 11778 37492 11788
rect 37548 11732 37604 12348
rect 37548 11666 37604 11676
rect 37660 12180 37716 12190
rect 37324 11508 37380 11518
rect 37660 11508 37716 12124
rect 37324 10388 37380 11452
rect 37548 11452 37716 11508
rect 37772 11508 37828 11518
rect 37436 11172 37492 11182
rect 37436 11078 37492 11116
rect 37548 11060 37604 11452
rect 37772 11394 37828 11452
rect 37772 11342 37774 11394
rect 37826 11342 37828 11394
rect 37772 11330 37828 11342
rect 37660 11284 37716 11294
rect 37660 11190 37716 11228
rect 37884 11284 37940 12460
rect 38108 12180 38164 12796
rect 38220 12404 38276 12414
rect 38332 12404 38388 12908
rect 38556 12898 38612 12908
rect 38668 12964 38724 12974
rect 38668 12870 38724 12908
rect 38780 12740 38836 12750
rect 38220 12402 38388 12404
rect 38220 12350 38222 12402
rect 38274 12350 38388 12402
rect 38220 12348 38388 12350
rect 38444 12404 38500 12414
rect 38220 12338 38276 12348
rect 38444 12310 38500 12348
rect 38668 12292 38724 12302
rect 38668 12198 38724 12236
rect 38108 12124 38276 12180
rect 38108 11956 38164 11966
rect 38108 11862 38164 11900
rect 38220 11394 38276 12124
rect 38220 11342 38222 11394
rect 38274 11342 38276 11394
rect 38220 11330 38276 11342
rect 38556 12068 38612 12078
rect 37884 11218 37940 11228
rect 38444 11284 38500 11322
rect 38444 11218 38500 11228
rect 38556 11282 38612 12012
rect 38780 12068 38836 12684
rect 38780 12002 38836 12012
rect 38892 11620 38948 13020
rect 39004 12852 39060 12862
rect 39004 12758 39060 12796
rect 38892 11564 39060 11620
rect 38556 11230 38558 11282
rect 38610 11230 38612 11282
rect 38444 11060 38500 11070
rect 38556 11060 38612 11230
rect 37548 11004 37716 11060
rect 37660 10836 37716 11004
rect 38500 11004 38612 11060
rect 38668 11508 38724 11518
rect 38332 10836 38388 10846
rect 37548 10780 37716 10836
rect 38220 10834 38388 10836
rect 38220 10782 38334 10834
rect 38386 10782 38388 10834
rect 38220 10780 38388 10782
rect 37436 10612 37492 10622
rect 37436 10518 37492 10556
rect 37324 10332 37492 10388
rect 37436 9604 37492 10332
rect 37548 10052 37604 10780
rect 37660 10612 37716 10622
rect 38108 10612 38164 10622
rect 37660 10518 37716 10556
rect 37772 10610 38164 10612
rect 37772 10558 38110 10610
rect 38162 10558 38164 10610
rect 37772 10556 38164 10558
rect 37660 10052 37716 10062
rect 37548 10050 37716 10052
rect 37548 9998 37662 10050
rect 37714 9998 37716 10050
rect 37548 9996 37716 9998
rect 37660 9986 37716 9996
rect 37772 10052 37828 10556
rect 38108 10546 38164 10556
rect 38220 10500 38276 10780
rect 38332 10770 38388 10780
rect 38444 10836 38500 11004
rect 38668 10836 38724 11452
rect 38444 10770 38500 10780
rect 38556 10780 38724 10836
rect 38892 11060 38948 11070
rect 38444 10612 38500 10622
rect 38220 10434 38276 10444
rect 38332 10610 38500 10612
rect 38332 10558 38446 10610
rect 38498 10558 38500 10610
rect 38332 10556 38500 10558
rect 37548 9828 37604 9838
rect 37548 9734 37604 9772
rect 37772 9826 37828 9996
rect 37772 9774 37774 9826
rect 37826 9774 37828 9826
rect 37772 9762 37828 9774
rect 37884 9940 37940 9950
rect 37436 9548 37604 9604
rect 37324 9492 37380 9502
rect 37324 9266 37380 9436
rect 37324 9214 37326 9266
rect 37378 9214 37380 9266
rect 37324 9202 37380 9214
rect 37436 9042 37492 9054
rect 37436 8990 37438 9042
rect 37490 8990 37492 9042
rect 37324 8820 37380 8830
rect 37324 8726 37380 8764
rect 37436 8484 37492 8990
rect 37324 8428 37492 8484
rect 37324 7812 37380 8428
rect 37436 8260 37492 8270
rect 37548 8260 37604 9548
rect 37436 8258 37604 8260
rect 37436 8206 37438 8258
rect 37490 8206 37604 8258
rect 37436 8204 37604 8206
rect 37660 9492 37716 9502
rect 37884 9492 37940 9884
rect 38332 9828 38388 10556
rect 38444 10546 38500 10556
rect 38556 10388 38612 10780
rect 37996 9772 38388 9828
rect 37996 9714 38052 9772
rect 37996 9662 37998 9714
rect 38050 9662 38052 9714
rect 37996 9650 38052 9662
rect 37884 9436 38164 9492
rect 37660 8708 37716 9436
rect 38108 9266 38164 9436
rect 38108 9214 38110 9266
rect 38162 9214 38164 9266
rect 38108 9202 38164 9214
rect 37996 9044 38052 9054
rect 37996 8950 38052 8988
rect 37436 8194 37492 8204
rect 37660 8146 37716 8652
rect 38108 8818 38164 8830
rect 38108 8766 38110 8818
rect 38162 8766 38164 8818
rect 38108 8708 38164 8766
rect 38108 8642 38164 8652
rect 38332 8484 38388 9772
rect 38444 10332 38612 10388
rect 38668 10610 38724 10622
rect 38668 10558 38670 10610
rect 38722 10558 38724 10610
rect 38444 8708 38500 10332
rect 38556 9828 38612 9838
rect 38668 9828 38724 10558
rect 38612 9772 38724 9828
rect 38780 9938 38836 9950
rect 38780 9886 38782 9938
rect 38834 9886 38836 9938
rect 38780 9828 38836 9886
rect 38556 9734 38612 9772
rect 38780 9762 38836 9772
rect 38444 8642 38500 8652
rect 38780 9602 38836 9614
rect 38780 9550 38782 9602
rect 38834 9550 38836 9602
rect 38444 8484 38500 8494
rect 37996 8482 38500 8484
rect 37996 8430 38446 8482
rect 38498 8430 38500 8482
rect 37996 8428 38500 8430
rect 37660 8094 37662 8146
rect 37714 8094 37716 8146
rect 37660 8082 37716 8094
rect 37772 8148 37828 8158
rect 37772 8054 37828 8092
rect 37324 7746 37380 7756
rect 37884 8036 37940 8046
rect 37884 7698 37940 7980
rect 37884 7646 37886 7698
rect 37938 7646 37940 7698
rect 37884 7634 37940 7646
rect 37996 7698 38052 8428
rect 38444 8418 38500 8428
rect 38668 8484 38724 8494
rect 37996 7646 37998 7698
rect 38050 7646 38052 7698
rect 37996 7634 38052 7646
rect 38108 8260 38164 8270
rect 38332 8260 38388 8270
rect 37212 7532 37828 7588
rect 37772 7476 37828 7532
rect 37772 7420 37940 7476
rect 37436 7364 37492 7374
rect 37100 7362 37492 7364
rect 37100 7310 37438 7362
rect 37490 7310 37492 7362
rect 37100 7308 37492 7310
rect 37436 7298 37492 7308
rect 37212 7140 37268 7150
rect 37212 6132 37268 7084
rect 37884 6578 37940 7420
rect 38108 6692 38164 8204
rect 37884 6526 37886 6578
rect 37938 6526 37940 6578
rect 37884 6514 37940 6526
rect 37996 6636 38164 6692
rect 38220 8204 38332 8260
rect 38220 7698 38276 8204
rect 38332 8194 38388 8204
rect 38220 7646 38222 7698
rect 38274 7646 38276 7698
rect 37772 6468 37828 6478
rect 37212 6066 37268 6076
rect 37324 6466 37828 6468
rect 37324 6414 37774 6466
rect 37826 6414 37828 6466
rect 37324 6412 37828 6414
rect 37324 6130 37380 6412
rect 37772 6402 37828 6412
rect 37996 6244 38052 6636
rect 38108 6468 38164 6478
rect 38220 6468 38276 7646
rect 38108 6466 38276 6468
rect 38108 6414 38110 6466
rect 38162 6414 38276 6466
rect 38108 6412 38276 6414
rect 38332 7812 38388 7822
rect 38108 6402 38164 6412
rect 37324 6078 37326 6130
rect 37378 6078 37380 6130
rect 37324 6066 37380 6078
rect 37548 6188 38052 6244
rect 37548 6130 37604 6188
rect 37548 6078 37550 6130
rect 37602 6078 37604 6130
rect 37548 6066 37604 6078
rect 38220 6132 38276 6142
rect 38220 6038 38276 6076
rect 37772 6020 37828 6030
rect 37772 5926 37828 5964
rect 37212 5906 37268 5918
rect 37212 5854 37214 5906
rect 37266 5854 37268 5906
rect 36988 3668 37044 5068
rect 37100 5236 37156 5246
rect 37100 4226 37156 5180
rect 37100 4174 37102 4226
rect 37154 4174 37156 4226
rect 37100 4162 37156 4174
rect 37100 3668 37156 3678
rect 36988 3666 37156 3668
rect 36988 3614 37102 3666
rect 37154 3614 37156 3666
rect 36988 3612 37156 3614
rect 37100 3602 37156 3612
rect 37212 3332 37268 5854
rect 37436 5796 37492 5806
rect 37436 5702 37492 5740
rect 37772 5796 37828 5806
rect 37660 5348 37716 5358
rect 37660 5234 37716 5292
rect 37660 5182 37662 5234
rect 37714 5182 37716 5234
rect 37660 5170 37716 5182
rect 37212 3266 37268 3276
rect 37436 4788 37492 4798
rect 36540 3042 36596 3052
rect 35420 2818 35476 2828
rect 35308 2594 35364 2604
rect 34748 800 34804 2380
rect 36092 2100 36148 2110
rect 36092 800 36148 2044
rect 37436 800 37492 4732
rect 37772 3780 37828 5740
rect 37772 3714 37828 3724
rect 38332 4676 38388 7756
rect 38556 7474 38612 7486
rect 38556 7422 38558 7474
rect 38610 7422 38612 7474
rect 38444 6692 38500 6702
rect 38444 6598 38500 6636
rect 38556 5348 38612 7422
rect 38556 5282 38612 5292
rect 38668 5236 38724 8428
rect 38780 8258 38836 9550
rect 38892 9266 38948 11004
rect 39004 9492 39060 11564
rect 39116 11284 39172 13020
rect 39340 12962 39396 13356
rect 39340 12910 39342 12962
rect 39394 12910 39396 12962
rect 39340 12898 39396 12910
rect 39452 12740 39508 13692
rect 39676 12964 39732 13804
rect 39676 12832 39732 12908
rect 40012 13412 40068 13422
rect 40012 12962 40068 13356
rect 40012 12910 40014 12962
rect 40066 12910 40068 12962
rect 39900 12852 39956 12862
rect 39900 12758 39956 12796
rect 39788 12740 39844 12750
rect 39452 12684 39732 12740
rect 39452 12404 39508 12414
rect 39452 12290 39508 12348
rect 39452 12238 39454 12290
rect 39506 12238 39508 12290
rect 39452 11788 39508 12238
rect 39116 11218 39172 11228
rect 39228 11732 39508 11788
rect 39676 12402 39732 12684
rect 39676 12350 39678 12402
rect 39730 12350 39732 12402
rect 39228 10834 39284 11732
rect 39452 11506 39508 11518
rect 39452 11454 39454 11506
rect 39506 11454 39508 11506
rect 39452 11396 39508 11454
rect 39452 11330 39508 11340
rect 39564 11170 39620 11182
rect 39564 11118 39566 11170
rect 39618 11118 39620 11170
rect 39564 10836 39620 11118
rect 39228 10782 39230 10834
rect 39282 10782 39284 10834
rect 39228 10770 39284 10782
rect 39452 10780 39564 10836
rect 39340 10722 39396 10734
rect 39340 10670 39342 10722
rect 39394 10670 39396 10722
rect 39004 9426 39060 9436
rect 39228 9492 39284 9502
rect 38892 9214 38894 9266
rect 38946 9214 38948 9266
rect 38892 9202 38948 9214
rect 39228 9268 39284 9436
rect 39228 9202 39284 9212
rect 39004 9042 39060 9054
rect 39004 8990 39006 9042
rect 39058 8990 39060 9042
rect 38780 8206 38782 8258
rect 38834 8206 38836 8258
rect 38780 6468 38836 8206
rect 38892 8818 38948 8830
rect 38892 8766 38894 8818
rect 38946 8766 38948 8818
rect 38892 7812 38948 8766
rect 39004 8484 39060 8990
rect 39340 8820 39396 10670
rect 39452 9492 39508 10780
rect 39564 10770 39620 10780
rect 39564 10610 39620 10622
rect 39564 10558 39566 10610
rect 39618 10558 39620 10610
rect 39564 9940 39620 10558
rect 39564 9874 39620 9884
rect 39676 9938 39732 12350
rect 39788 12066 39844 12684
rect 39788 12014 39790 12066
rect 39842 12014 39844 12066
rect 39788 12002 39844 12014
rect 40012 11620 40068 12910
rect 40012 11554 40068 11564
rect 39788 11396 39844 11434
rect 39788 11330 39844 11340
rect 39788 10610 39844 10622
rect 39788 10558 39790 10610
rect 39842 10558 39844 10610
rect 39788 10164 39844 10558
rect 39788 10098 39844 10108
rect 40124 9940 40180 17724
rect 40236 15540 40292 18732
rect 40348 18226 40404 18844
rect 40460 18564 40516 18956
rect 40740 18956 40852 19012
rect 41020 19010 41300 19012
rect 41020 18958 41246 19010
rect 41298 18958 41300 19010
rect 41020 18956 41300 18958
rect 40684 18918 40740 18956
rect 40460 18498 40516 18508
rect 40684 18452 40740 18462
rect 40348 18174 40350 18226
rect 40402 18174 40404 18226
rect 40348 18162 40404 18174
rect 40460 18338 40516 18350
rect 40460 18286 40462 18338
rect 40514 18286 40516 18338
rect 40460 17892 40516 18286
rect 40460 17332 40516 17836
rect 40460 17266 40516 17276
rect 40572 17554 40628 17566
rect 40572 17502 40574 17554
rect 40626 17502 40628 17554
rect 40572 17220 40628 17502
rect 40572 17154 40628 17164
rect 40684 17442 40740 18396
rect 40796 18340 40852 18350
rect 40796 18226 40852 18284
rect 40796 18174 40798 18226
rect 40850 18174 40852 18226
rect 40796 18162 40852 18174
rect 40684 17390 40686 17442
rect 40738 17390 40740 17442
rect 40572 16996 40628 17006
rect 40572 16902 40628 16940
rect 40460 16884 40516 16894
rect 40460 16790 40516 16828
rect 40348 16548 40404 16558
rect 40348 15764 40404 16492
rect 40572 15988 40628 16026
rect 40572 15922 40628 15932
rect 40348 15698 40404 15708
rect 40460 15874 40516 15886
rect 40460 15822 40462 15874
rect 40514 15822 40516 15874
rect 40460 15652 40516 15822
rect 40460 15586 40516 15596
rect 40572 15764 40628 15774
rect 40236 15474 40292 15484
rect 40572 15538 40628 15708
rect 40572 15486 40574 15538
rect 40626 15486 40628 15538
rect 40572 15474 40628 15486
rect 40348 15426 40404 15438
rect 40348 15374 40350 15426
rect 40402 15374 40404 15426
rect 40236 15316 40292 15326
rect 40236 15222 40292 15260
rect 40236 14644 40292 14654
rect 40236 11508 40292 14588
rect 40348 14530 40404 15374
rect 40684 15316 40740 17390
rect 41020 16660 41076 18956
rect 41244 18946 41300 18956
rect 41356 18228 41412 19180
rect 41020 16594 41076 16604
rect 41132 18172 41412 18228
rect 41020 15876 41076 15886
rect 41020 15782 41076 15820
rect 40684 15250 40740 15260
rect 40348 14478 40350 14530
rect 40402 14478 40404 14530
rect 40348 14466 40404 14478
rect 40684 14420 40740 14430
rect 40740 14364 40852 14420
rect 40572 14306 40628 14318
rect 40572 14254 40574 14306
rect 40626 14254 40628 14306
rect 40684 14288 40740 14364
rect 40572 13972 40628 14254
rect 40572 13906 40628 13916
rect 40684 14196 40740 14206
rect 40684 13858 40740 14140
rect 40684 13806 40686 13858
rect 40738 13806 40740 13858
rect 40572 13748 40628 13758
rect 40572 13654 40628 13692
rect 40684 13636 40740 13806
rect 40684 13570 40740 13580
rect 40572 12964 40628 12974
rect 40572 12870 40628 12908
rect 40684 12740 40740 12750
rect 40684 12646 40740 12684
rect 40572 12628 40628 12638
rect 40460 12290 40516 12302
rect 40460 12238 40462 12290
rect 40514 12238 40516 12290
rect 40460 12180 40516 12238
rect 40572 12290 40628 12572
rect 40572 12238 40574 12290
rect 40626 12238 40628 12290
rect 40572 12226 40628 12238
rect 40460 12114 40516 12124
rect 40460 11956 40516 11966
rect 40236 11442 40292 11452
rect 40348 11954 40516 11956
rect 40348 11902 40462 11954
rect 40514 11902 40516 11954
rect 40348 11900 40516 11902
rect 40236 11060 40292 11070
rect 40236 10834 40292 11004
rect 40348 10948 40404 11900
rect 40460 11890 40516 11900
rect 40460 11620 40516 11630
rect 40460 11526 40516 11564
rect 40460 11284 40516 11294
rect 40460 11190 40516 11228
rect 40572 11282 40628 11294
rect 40572 11230 40574 11282
rect 40626 11230 40628 11282
rect 40572 11172 40628 11230
rect 40572 11106 40628 11116
rect 40796 10948 40852 14364
rect 40908 13748 40964 13758
rect 40908 13746 41076 13748
rect 40908 13694 40910 13746
rect 40962 13694 41076 13746
rect 40908 13692 41076 13694
rect 40908 13682 40964 13692
rect 40908 12738 40964 12750
rect 40908 12686 40910 12738
rect 40962 12686 40964 12738
rect 40908 12292 40964 12686
rect 41020 12404 41076 13692
rect 41020 12338 41076 12348
rect 40908 12226 40964 12236
rect 40348 10882 40404 10892
rect 40460 10892 40852 10948
rect 41020 11172 41076 11182
rect 41132 11172 41188 18172
rect 41244 18004 41300 18014
rect 41244 17890 41300 17948
rect 41244 17838 41246 17890
rect 41298 17838 41300 17890
rect 41244 17826 41300 17838
rect 41356 17778 41412 18172
rect 41356 17726 41358 17778
rect 41410 17726 41412 17778
rect 41356 17714 41412 17726
rect 41468 18340 41524 18350
rect 41356 17444 41412 17454
rect 41244 17108 41300 17118
rect 41244 13748 41300 17052
rect 41356 14308 41412 17388
rect 41468 16100 41524 18284
rect 41580 17780 41636 20860
rect 41916 19908 41972 21420
rect 42028 20916 42084 20926
rect 42028 20822 42084 20860
rect 41804 19906 41972 19908
rect 41804 19854 41918 19906
rect 41970 19854 41972 19906
rect 41804 19852 41972 19854
rect 41692 19010 41748 19022
rect 41692 18958 41694 19010
rect 41746 18958 41748 19010
rect 41692 17892 41748 18958
rect 41804 18228 41860 19852
rect 41916 19842 41972 19852
rect 41804 18162 41860 18172
rect 41916 19458 41972 19470
rect 41916 19406 41918 19458
rect 41970 19406 41972 19458
rect 41916 18450 41972 19406
rect 42028 19348 42084 19358
rect 42028 19254 42084 19292
rect 41916 18398 41918 18450
rect 41970 18398 41972 18450
rect 41916 18116 41972 18398
rect 42028 18340 42084 18350
rect 42028 18246 42084 18284
rect 41916 18050 41972 18060
rect 41692 17826 41748 17836
rect 41916 17892 41972 17902
rect 41580 17714 41636 17724
rect 41916 17778 41972 17836
rect 42028 17892 42084 17902
rect 42140 17892 42196 21756
rect 42028 17890 42196 17892
rect 42028 17838 42030 17890
rect 42082 17838 42196 17890
rect 42028 17836 42196 17838
rect 42028 17826 42084 17836
rect 41916 17726 41918 17778
rect 41970 17726 41972 17778
rect 41916 17714 41972 17726
rect 41916 17332 41972 17342
rect 41468 16034 41524 16044
rect 41580 17220 41636 17230
rect 41580 15988 41636 17164
rect 41804 16996 41860 17006
rect 41692 16994 41860 16996
rect 41692 16942 41806 16994
rect 41858 16942 41860 16994
rect 41692 16940 41860 16942
rect 41692 16660 41748 16940
rect 41804 16930 41860 16940
rect 41916 16994 41972 17276
rect 41916 16942 41918 16994
rect 41970 16942 41972 16994
rect 41916 16930 41972 16942
rect 41692 16594 41748 16604
rect 41804 16772 41860 16782
rect 41804 16658 41860 16716
rect 41804 16606 41806 16658
rect 41858 16606 41860 16658
rect 41804 16594 41860 16606
rect 41916 16436 41972 16446
rect 41804 16100 41860 16110
rect 41804 16006 41860 16044
rect 41692 15988 41748 15998
rect 41580 15986 41748 15988
rect 41580 15934 41694 15986
rect 41746 15934 41748 15986
rect 41580 15932 41748 15934
rect 41468 15876 41524 15886
rect 41468 15782 41524 15820
rect 41580 15540 41636 15932
rect 41692 15922 41748 15932
rect 41468 15484 41636 15540
rect 41804 15540 41860 15550
rect 41916 15540 41972 16380
rect 41804 15538 41972 15540
rect 41804 15486 41806 15538
rect 41858 15486 41972 15538
rect 41804 15484 41972 15486
rect 41468 15204 41524 15484
rect 41804 15474 41860 15484
rect 41692 15370 41748 15382
rect 41692 15318 41694 15370
rect 41746 15318 41748 15370
rect 41692 15316 41748 15318
rect 41692 15204 41748 15260
rect 41468 15138 41524 15148
rect 41580 15148 41748 15204
rect 41804 15204 41860 15214
rect 41356 14242 41412 14252
rect 41468 14306 41524 14318
rect 41468 14254 41470 14306
rect 41522 14254 41524 14306
rect 41468 13748 41524 14254
rect 41580 14196 41636 15148
rect 41804 14530 41860 15148
rect 41804 14478 41806 14530
rect 41858 14478 41860 14530
rect 41804 14466 41860 14478
rect 41916 14532 41972 15484
rect 41916 14466 41972 14476
rect 42028 15874 42084 15886
rect 42028 15822 42030 15874
rect 42082 15822 42084 15874
rect 42028 15538 42084 15822
rect 42028 15486 42030 15538
rect 42082 15486 42084 15538
rect 41692 14308 41748 14318
rect 41748 14252 41972 14308
rect 41692 14176 41748 14252
rect 41580 14130 41636 14140
rect 41692 13972 41748 13982
rect 41748 13916 41860 13972
rect 41692 13878 41748 13916
rect 41580 13748 41636 13758
rect 41244 13682 41300 13692
rect 41356 13746 41636 13748
rect 41356 13694 41582 13746
rect 41634 13694 41636 13746
rect 41356 13692 41636 13694
rect 41356 11394 41412 13692
rect 41580 13682 41636 13692
rect 41692 13524 41748 13534
rect 41580 13522 41748 13524
rect 41580 13470 41694 13522
rect 41746 13470 41748 13522
rect 41580 13468 41748 13470
rect 41468 12964 41524 12974
rect 41468 12870 41524 12908
rect 41356 11342 41358 11394
rect 41410 11342 41412 11394
rect 41356 11330 41412 11342
rect 41244 11284 41300 11294
rect 41244 11190 41300 11228
rect 41020 11170 41188 11172
rect 41020 11118 41022 11170
rect 41074 11118 41188 11170
rect 41020 11116 41188 11118
rect 40236 10782 40238 10834
rect 40290 10782 40292 10834
rect 40236 10770 40292 10782
rect 40348 10724 40404 10734
rect 40460 10724 40516 10892
rect 40348 10722 40516 10724
rect 40348 10670 40350 10722
rect 40402 10670 40516 10722
rect 40348 10668 40516 10670
rect 40348 10658 40404 10668
rect 40572 10612 40628 10622
rect 40572 10610 40740 10612
rect 40572 10558 40574 10610
rect 40626 10558 40740 10610
rect 40572 10556 40740 10558
rect 40572 10546 40628 10556
rect 40460 10500 40516 10510
rect 39676 9886 39678 9938
rect 39730 9886 39732 9938
rect 39676 9874 39732 9886
rect 40012 9884 40180 9940
rect 40348 10052 40404 10062
rect 39788 9826 39844 9838
rect 39788 9774 39790 9826
rect 39842 9774 39844 9826
rect 39564 9716 39620 9726
rect 39564 9714 39732 9716
rect 39564 9662 39566 9714
rect 39618 9662 39732 9714
rect 39564 9660 39732 9662
rect 39564 9650 39620 9660
rect 39676 9492 39732 9660
rect 39788 9604 39844 9774
rect 39788 9538 39844 9548
rect 39452 9436 39620 9492
rect 39452 9268 39508 9278
rect 39452 9174 39508 9212
rect 39340 8754 39396 8764
rect 39004 8418 39060 8428
rect 39340 8596 39396 8606
rect 39004 8146 39060 8158
rect 39004 8094 39006 8146
rect 39058 8094 39060 8146
rect 39004 8036 39060 8094
rect 39004 7970 39060 7980
rect 38892 7746 38948 7756
rect 39116 7700 39172 7710
rect 39116 7606 39172 7644
rect 39340 7586 39396 8540
rect 39564 8372 39620 9436
rect 39676 9426 39732 9436
rect 39900 9492 39956 9502
rect 39788 9380 39844 9390
rect 39676 9154 39732 9166
rect 39676 9102 39678 9154
rect 39730 9102 39732 9154
rect 39676 9044 39732 9102
rect 39788 9154 39844 9324
rect 39788 9102 39790 9154
rect 39842 9102 39844 9154
rect 39788 9090 39844 9102
rect 39676 8978 39732 8988
rect 39564 8306 39620 8316
rect 39340 7534 39342 7586
rect 39394 7534 39396 7586
rect 39340 7522 39396 7534
rect 39452 8258 39508 8270
rect 39788 8260 39844 8270
rect 39452 8206 39454 8258
rect 39506 8206 39508 8258
rect 39228 7364 39284 7374
rect 39452 7364 39508 8206
rect 39676 8258 39844 8260
rect 39676 8206 39790 8258
rect 39842 8206 39844 8258
rect 39676 8204 39844 8206
rect 39676 8148 39732 8204
rect 39788 8194 39844 8204
rect 39676 8082 39732 8092
rect 39228 7362 39508 7364
rect 39228 7310 39230 7362
rect 39282 7310 39508 7362
rect 39228 7308 39508 7310
rect 39788 8036 39844 8046
rect 39228 6916 39284 7308
rect 39228 6850 39284 6860
rect 38780 6402 38836 6412
rect 39004 6802 39060 6814
rect 39004 6750 39006 6802
rect 39058 6750 39060 6802
rect 38892 5796 38948 5806
rect 38892 5702 38948 5740
rect 38668 5180 38836 5236
rect 38780 4788 38836 5180
rect 38332 3556 38388 4620
rect 38668 4732 38836 4788
rect 38892 5010 38948 5022
rect 38892 4958 38894 5010
rect 38946 4958 38948 5010
rect 38892 4788 38948 4958
rect 38332 3490 38388 3500
rect 38444 4450 38500 4462
rect 38444 4398 38446 4450
rect 38498 4398 38500 4450
rect 38108 3444 38164 3482
rect 38108 3378 38164 3388
rect 38444 2884 38500 4398
rect 38444 2100 38500 2828
rect 38444 2034 38500 2044
rect 38668 1652 38724 4732
rect 38892 4722 38948 4732
rect 38668 1586 38724 1596
rect 38780 4452 38836 4462
rect 38780 2996 38836 4396
rect 39004 3780 39060 6750
rect 39116 5460 39172 5470
rect 39116 4226 39172 5404
rect 39116 4174 39118 4226
rect 39170 4174 39172 4226
rect 39116 4162 39172 4174
rect 39676 5234 39732 5246
rect 39676 5182 39678 5234
rect 39730 5182 39732 5234
rect 39676 4228 39732 5182
rect 39788 5012 39844 7980
rect 39900 7700 39956 9436
rect 39900 7586 39956 7644
rect 40012 7698 40068 9884
rect 40348 9828 40404 9996
rect 40124 9716 40180 9726
rect 40124 9714 40292 9716
rect 40124 9662 40126 9714
rect 40178 9662 40292 9714
rect 40124 9660 40292 9662
rect 40124 9650 40180 9660
rect 40124 8146 40180 8158
rect 40124 8094 40126 8146
rect 40178 8094 40180 8146
rect 40124 7812 40180 8094
rect 40236 8036 40292 9660
rect 40348 8708 40404 9772
rect 40460 9266 40516 10444
rect 40572 9716 40628 9726
rect 40572 9622 40628 9660
rect 40460 9214 40462 9266
rect 40514 9214 40516 9266
rect 40460 9202 40516 9214
rect 40572 9156 40628 9166
rect 40572 9062 40628 9100
rect 40460 9044 40516 9054
rect 40460 8818 40516 8988
rect 40684 8932 40740 10556
rect 40796 10610 40852 10622
rect 40796 10558 40798 10610
rect 40850 10558 40852 10610
rect 40796 10052 40852 10558
rect 40796 9986 40852 9996
rect 40908 10164 40964 10174
rect 40796 9828 40852 9838
rect 40796 9714 40852 9772
rect 40908 9826 40964 10108
rect 40908 9774 40910 9826
rect 40962 9774 40964 9826
rect 40908 9762 40964 9774
rect 40796 9662 40798 9714
rect 40850 9662 40852 9714
rect 40796 9044 40852 9662
rect 40796 8978 40852 8988
rect 40908 9604 40964 9614
rect 40460 8766 40462 8818
rect 40514 8766 40516 8818
rect 40460 8754 40516 8766
rect 40572 8876 40740 8932
rect 40348 8642 40404 8652
rect 40236 7970 40292 7980
rect 40348 8372 40404 8382
rect 40124 7746 40180 7756
rect 40012 7646 40014 7698
rect 40066 7646 40068 7698
rect 40012 7634 40068 7646
rect 39900 7534 39902 7586
rect 39954 7534 39956 7586
rect 39900 7522 39956 7534
rect 40236 7476 40292 7486
rect 40348 7476 40404 8316
rect 40236 7474 40404 7476
rect 40236 7422 40238 7474
rect 40290 7422 40404 7474
rect 40236 7420 40404 7422
rect 40236 7410 40292 7420
rect 40572 6916 40628 8876
rect 40684 8372 40740 8382
rect 40684 8278 40740 8316
rect 40684 7476 40740 7486
rect 40684 7362 40740 7420
rect 40684 7310 40686 7362
rect 40738 7310 40740 7362
rect 40684 7140 40740 7310
rect 40684 7074 40740 7084
rect 40572 6850 40628 6860
rect 40796 6804 40852 6814
rect 39900 6580 39956 6590
rect 39900 6486 39956 6524
rect 40796 6130 40852 6748
rect 40908 6690 40964 9548
rect 41020 8596 41076 11116
rect 41468 10052 41524 10062
rect 41356 9604 41412 9614
rect 41356 9510 41412 9548
rect 41468 9380 41524 9996
rect 41580 9940 41636 13468
rect 41692 13458 41748 13468
rect 41692 13300 41748 13310
rect 41692 12738 41748 13244
rect 41692 12686 41694 12738
rect 41746 12686 41748 12738
rect 41692 12628 41748 12686
rect 41692 12562 41748 12572
rect 41804 12962 41860 13916
rect 41916 13412 41972 14252
rect 41916 13346 41972 13356
rect 41804 12910 41806 12962
rect 41858 12910 41860 12962
rect 41692 12404 41748 12414
rect 41692 12310 41748 12348
rect 41804 12290 41860 12910
rect 42028 12964 42084 15486
rect 42140 13300 42196 17836
rect 42252 21924 42308 21934
rect 42252 17668 42308 21868
rect 42364 20916 42420 23212
rect 42364 20850 42420 20860
rect 42476 18004 42532 24108
rect 42812 23940 42868 23950
rect 42476 17938 42532 17948
rect 42588 22372 42644 22382
rect 42252 15874 42308 17612
rect 42252 15822 42254 15874
rect 42306 15822 42308 15874
rect 42252 15810 42308 15822
rect 42140 13234 42196 13244
rect 42364 14084 42420 14094
rect 42252 13076 42308 13086
rect 42028 12908 42196 12964
rect 41804 12238 41806 12290
rect 41858 12238 41860 12290
rect 41804 12226 41860 12238
rect 42028 12740 42084 12750
rect 41916 12068 41972 12078
rect 41692 11956 41748 11966
rect 41692 11954 41860 11956
rect 41692 11902 41694 11954
rect 41746 11902 41860 11954
rect 41692 11900 41860 11902
rect 41692 11890 41748 11900
rect 41692 10836 41748 10846
rect 41692 10742 41748 10780
rect 41804 10724 41860 11900
rect 41916 11618 41972 12012
rect 41916 11566 41918 11618
rect 41970 11566 41972 11618
rect 41916 11554 41972 11566
rect 42028 11506 42084 12684
rect 42028 11454 42030 11506
rect 42082 11454 42084 11506
rect 42028 11442 42084 11454
rect 42140 11284 42196 12908
rect 42140 11218 42196 11228
rect 41804 10722 41972 10724
rect 41804 10670 41806 10722
rect 41858 10670 41972 10722
rect 41804 10668 41972 10670
rect 41804 10658 41860 10668
rect 41692 10388 41748 10398
rect 41692 10294 41748 10332
rect 41580 9884 41860 9940
rect 41692 9716 41748 9726
rect 41692 9622 41748 9660
rect 41580 9602 41636 9614
rect 41580 9550 41582 9602
rect 41634 9550 41636 9602
rect 41580 9492 41636 9550
rect 41804 9604 41860 9884
rect 41916 9828 41972 10668
rect 41916 9762 41972 9772
rect 41804 9548 42084 9604
rect 41580 9436 41972 9492
rect 41468 9324 41636 9380
rect 41468 9044 41524 9054
rect 41020 8530 41076 8540
rect 41132 9042 41524 9044
rect 41132 8990 41470 9042
rect 41522 8990 41524 9042
rect 41132 8988 41524 8990
rect 41020 8148 41076 8158
rect 41020 8054 41076 8092
rect 40908 6638 40910 6690
rect 40962 6638 40964 6690
rect 40908 6626 40964 6638
rect 41020 6580 41076 6590
rect 41132 6580 41188 8988
rect 41468 8978 41524 8988
rect 41356 8820 41412 8830
rect 41244 8708 41300 8718
rect 41244 7700 41300 8652
rect 41244 7634 41300 7644
rect 41356 7252 41412 8764
rect 41580 8484 41636 9324
rect 41804 9268 41860 9278
rect 41692 9156 41748 9166
rect 41692 9062 41748 9100
rect 41804 9154 41860 9212
rect 41804 9102 41806 9154
rect 41858 9102 41860 9154
rect 41804 9090 41860 9102
rect 41692 8484 41748 8494
rect 41580 8482 41748 8484
rect 41580 8430 41694 8482
rect 41746 8430 41748 8482
rect 41580 8428 41748 8430
rect 41692 8418 41748 8428
rect 41356 7186 41412 7196
rect 41468 8148 41524 8158
rect 41020 6578 41188 6580
rect 41020 6526 41022 6578
rect 41074 6526 41188 6578
rect 41020 6524 41188 6526
rect 41020 6514 41076 6524
rect 40796 6078 40798 6130
rect 40850 6078 40852 6130
rect 40796 6066 40852 6078
rect 41244 6468 41300 6478
rect 40124 6020 40180 6030
rect 40124 5926 40180 5964
rect 41132 6020 41188 6030
rect 39788 4946 39844 4956
rect 40684 5010 40740 5022
rect 40684 4958 40686 5010
rect 40738 4958 40740 5010
rect 40236 4900 40292 4910
rect 40124 4452 40180 4462
rect 40124 4358 40180 4396
rect 39676 4162 39732 4172
rect 39004 3714 39060 3724
rect 39788 3780 39844 3790
rect 39116 3556 39172 3566
rect 39116 3462 39172 3500
rect 39564 3556 39620 3566
rect 39340 3444 39396 3482
rect 39564 3462 39620 3500
rect 39788 3554 39844 3724
rect 39788 3502 39790 3554
rect 39842 3502 39844 3554
rect 39788 3490 39844 3502
rect 39340 3378 39396 3388
rect 40124 3332 40180 3342
rect 40124 3238 40180 3276
rect 40236 3108 40292 4844
rect 40684 4900 40740 4958
rect 40684 4834 40740 4844
rect 40908 3556 40964 3566
rect 40908 3462 40964 3500
rect 41132 3388 41188 5964
rect 41244 5124 41300 6412
rect 41468 6130 41524 8092
rect 41692 8148 41748 8158
rect 41692 8054 41748 8092
rect 41804 8148 41860 8158
rect 41916 8148 41972 9436
rect 41804 8146 41972 8148
rect 41804 8094 41806 8146
rect 41858 8094 41972 8146
rect 41804 8092 41972 8094
rect 41580 8036 41636 8046
rect 41580 6690 41636 7980
rect 41804 7924 41860 8092
rect 42028 8036 42084 9548
rect 41804 7858 41860 7868
rect 41916 7980 42084 8036
rect 42140 8932 42196 8942
rect 41916 7812 41972 7980
rect 41692 7700 41748 7710
rect 41692 7606 41748 7644
rect 41804 7588 41860 7598
rect 41916 7588 41972 7756
rect 41804 7586 41972 7588
rect 41804 7534 41806 7586
rect 41858 7534 41972 7586
rect 41804 7532 41972 7534
rect 41804 7522 41860 7532
rect 41916 7364 41972 7374
rect 41692 7252 41748 7262
rect 41692 7158 41748 7196
rect 41580 6638 41582 6690
rect 41634 6638 41636 6690
rect 41580 6626 41636 6638
rect 41804 6916 41860 6926
rect 41804 6578 41860 6860
rect 41916 6690 41972 7308
rect 41916 6638 41918 6690
rect 41970 6638 41972 6690
rect 41916 6626 41972 6638
rect 42028 7140 42084 7150
rect 41804 6526 41806 6578
rect 41858 6526 41860 6578
rect 41804 6514 41860 6526
rect 41804 6244 41860 6254
rect 41468 6078 41470 6130
rect 41522 6078 41524 6130
rect 41468 6066 41524 6078
rect 41692 6132 41748 6142
rect 41692 6038 41748 6076
rect 41804 6018 41860 6188
rect 41804 5966 41806 6018
rect 41858 5966 41860 6018
rect 41804 5954 41860 5966
rect 41804 5348 41860 5358
rect 41804 5254 41860 5292
rect 41244 5058 41300 5068
rect 41580 5236 41636 5246
rect 41580 4450 41636 5180
rect 41916 5124 41972 5134
rect 41916 5030 41972 5068
rect 41804 5012 41860 5022
rect 41804 4918 41860 4956
rect 41580 4398 41582 4450
rect 41634 4398 41636 4450
rect 41580 4386 41636 4398
rect 41804 4340 41860 4350
rect 41804 4246 41860 4284
rect 41580 3780 41636 3790
rect 41356 3556 41412 3566
rect 41356 3462 41412 3500
rect 41580 3554 41636 3724
rect 42028 3666 42084 7084
rect 42140 6132 42196 8876
rect 42140 6066 42196 6076
rect 42252 4564 42308 13020
rect 42252 4498 42308 4508
rect 42364 3780 42420 14028
rect 42588 13972 42644 22316
rect 42476 13916 42644 13972
rect 42700 22148 42756 22158
rect 42476 8484 42532 13916
rect 42476 8418 42532 8428
rect 42588 13748 42644 13758
rect 42364 3714 42420 3724
rect 42028 3614 42030 3666
rect 42082 3614 42084 3666
rect 42028 3602 42084 3614
rect 41580 3502 41582 3554
rect 41634 3502 41636 3554
rect 41580 3490 41636 3502
rect 41468 3442 41524 3454
rect 41468 3390 41470 3442
rect 41522 3390 41524 3442
rect 41132 3332 41300 3388
rect 38780 800 38836 2940
rect 40124 3052 40292 3108
rect 41244 3108 41300 3332
rect 41468 3332 41524 3390
rect 41468 3266 41524 3276
rect 41244 3052 41524 3108
rect 40124 800 40180 3052
rect 41468 800 41524 3052
rect 42588 2548 42644 13692
rect 42588 2482 42644 2492
rect 42700 1540 42756 22092
rect 42812 13076 42868 23884
rect 42812 13010 42868 13020
rect 42924 23828 42980 23838
rect 42700 1474 42756 1484
rect 42812 6580 42868 6590
rect 42812 800 42868 6524
rect 42924 4788 42980 23772
rect 42924 4722 42980 4732
rect 43036 23044 43092 23054
rect 43036 2884 43092 22988
rect 43148 16996 43204 24444
rect 43148 16930 43204 16940
rect 43260 10276 43316 25228
rect 43260 10210 43316 10220
rect 43372 16884 43428 16894
rect 43036 2818 43092 2828
rect 43372 2660 43428 16828
rect 43372 2594 43428 2604
rect 1120 0 1232 800
rect 2464 0 2576 800
rect 3808 0 3920 800
rect 5152 0 5264 800
rect 6496 0 6608 800
rect 7840 0 7952 800
rect 9184 0 9296 800
rect 10528 0 10640 800
rect 11872 0 11984 800
rect 13216 0 13328 800
rect 14560 0 14672 800
rect 15904 0 16016 800
rect 17248 0 17360 800
rect 18592 0 18704 800
rect 19936 0 20048 800
rect 21280 0 21392 800
rect 22624 0 22736 800
rect 23968 0 24080 800
rect 25312 0 25424 800
rect 26656 0 26768 800
rect 28000 0 28112 800
rect 29344 0 29456 800
rect 30688 0 30800 800
rect 32032 0 32144 800
rect 33376 0 33488 800
rect 34720 0 34832 800
rect 36064 0 36176 800
rect 37408 0 37520 800
rect 38752 0 38864 800
rect 40096 0 40208 800
rect 41440 0 41552 800
rect 42784 0 42896 800
<< via2 >>
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 18396 39004 18452 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14364 24780 14420 24836
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 3388 22316 3444 22372
rect 8428 22316 8484 22372
rect 1820 21980 1876 22036
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1596 20860 1652 20916
rect 1148 4172 1204 4228
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1596 2604 1652 2660
rect 1708 18284 1764 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6748 15820 6804 15876
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 6412 13804 6468 13860
rect 3948 13692 4004 13748
rect 2940 13580 2996 13636
rect 2044 12572 2100 12628
rect 1820 9436 1876 9492
rect 1932 9100 1988 9156
rect 1932 8258 1988 8260
rect 1932 8206 1934 8258
rect 1934 8206 1986 8258
rect 1986 8206 1988 8258
rect 1932 8204 1988 8206
rect 2828 11900 2884 11956
rect 2716 10834 2772 10836
rect 2716 10782 2718 10834
rect 2718 10782 2770 10834
rect 2770 10782 2772 10834
rect 2716 10780 2772 10782
rect 2604 9324 2660 9380
rect 2156 8316 2212 8372
rect 2044 6076 2100 6132
rect 2156 7980 2212 8036
rect 2268 7868 2324 7924
rect 2828 8034 2884 8036
rect 2828 7982 2830 8034
rect 2830 7982 2882 8034
rect 2882 7982 2884 8034
rect 2828 7980 2884 7982
rect 2492 7196 2548 7252
rect 2604 7756 2660 7812
rect 2716 7698 2772 7700
rect 2716 7646 2718 7698
rect 2718 7646 2770 7698
rect 2770 7646 2772 7698
rect 2716 7644 2772 7646
rect 2716 6188 2772 6244
rect 3612 11170 3668 11172
rect 3612 11118 3614 11170
rect 3614 11118 3666 11170
rect 3666 11118 3668 11170
rect 3612 11116 3668 11118
rect 3276 9996 3332 10052
rect 3612 9996 3668 10052
rect 3836 9772 3892 9828
rect 3612 9436 3668 9492
rect 3836 9548 3892 9604
rect 3052 8930 3108 8932
rect 3052 8878 3054 8930
rect 3054 8878 3106 8930
rect 3106 8878 3108 8930
rect 3052 8876 3108 8878
rect 3500 8764 3556 8820
rect 3164 8316 3220 8372
rect 3052 8204 3108 8260
rect 3164 6636 3220 6692
rect 3724 9100 3780 9156
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5964 13244 6020 13300
rect 11340 20636 11396 20692
rect 10108 15148 10164 15204
rect 8428 14924 8484 14980
rect 9660 15036 9716 15092
rect 9100 13804 9156 13860
rect 7196 13244 7252 13300
rect 4284 11900 4340 11956
rect 4060 11170 4116 11172
rect 4060 11118 4062 11170
rect 4062 11118 4114 11170
rect 4114 11118 4116 11170
rect 4060 11116 4116 11118
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4508 11170 4564 11172
rect 4508 11118 4510 11170
rect 4510 11118 4562 11170
rect 4562 11118 4564 11170
rect 4508 11116 4564 11118
rect 4956 11004 5012 11060
rect 5292 11116 5348 11172
rect 5180 10780 5236 10836
rect 4060 10498 4116 10500
rect 4060 10446 4062 10498
rect 4062 10446 4114 10498
rect 4114 10446 4116 10498
rect 4060 10444 4116 10446
rect 4284 10332 4340 10388
rect 4172 9602 4228 9604
rect 4172 9550 4174 9602
rect 4174 9550 4226 9602
rect 4226 9550 4228 9602
rect 4172 9548 4228 9550
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4508 9996 4564 10052
rect 4396 9324 4452 9380
rect 4060 8876 4116 8932
rect 4284 8930 4340 8932
rect 4284 8878 4286 8930
rect 4286 8878 4338 8930
rect 4338 8878 4340 8930
rect 4284 8876 4340 8878
rect 5068 9938 5124 9940
rect 5068 9886 5070 9938
rect 5070 9886 5122 9938
rect 5122 9886 5124 9938
rect 5068 9884 5124 9886
rect 4844 9660 4900 9716
rect 4844 9100 4900 9156
rect 4172 8258 4228 8260
rect 4172 8206 4174 8258
rect 4174 8206 4226 8258
rect 4226 8206 4228 8258
rect 4172 8204 4228 8206
rect 3612 7644 3668 7700
rect 3724 7586 3780 7588
rect 3724 7534 3726 7586
rect 3726 7534 3778 7586
rect 3778 7534 3780 7586
rect 3724 7532 3780 7534
rect 3612 6748 3668 6804
rect 3164 6130 3220 6132
rect 3164 6078 3166 6130
rect 3166 6078 3218 6130
rect 3218 6078 3220 6130
rect 3164 6076 3220 6078
rect 3164 5292 3220 5348
rect 2940 5180 2996 5236
rect 1820 4620 1876 4676
rect 1932 4226 1988 4228
rect 1932 4174 1934 4226
rect 1934 4174 1986 4226
rect 1986 4174 1988 4226
rect 1932 4172 1988 4174
rect 1708 2380 1764 2436
rect 3612 5068 3668 5124
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4732 8316 4788 8372
rect 4508 7756 4564 7812
rect 4396 7474 4452 7476
rect 4396 7422 4398 7474
rect 4398 7422 4450 7474
rect 4450 7422 4452 7474
rect 4396 7420 4452 7422
rect 5068 8540 5124 8596
rect 4844 8204 4900 8260
rect 4956 8428 5012 8484
rect 5068 8316 5124 8372
rect 5292 9212 5348 9268
rect 5404 9154 5460 9156
rect 5404 9102 5406 9154
rect 5406 9102 5458 9154
rect 5458 9102 5460 9154
rect 5404 9100 5460 9102
rect 5292 8428 5348 8484
rect 4620 7644 4676 7700
rect 5068 7756 5124 7812
rect 5180 7980 5236 8036
rect 5180 7308 5236 7364
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4844 7084 4900 7140
rect 4684 7028 4740 7030
rect 4844 6578 4900 6580
rect 4844 6526 4846 6578
rect 4846 6526 4898 6578
rect 4898 6526 4900 6578
rect 4844 6524 4900 6526
rect 4172 6412 4228 6468
rect 3836 5404 3892 5460
rect 3948 5852 4004 5908
rect 3948 5346 4004 5348
rect 3948 5294 3950 5346
rect 3950 5294 4002 5346
rect 4002 5294 4004 5346
rect 3948 5292 4004 5294
rect 4060 5516 4116 5572
rect 3724 4284 3780 4340
rect 4060 4732 4116 4788
rect 3948 4450 4004 4452
rect 3948 4398 3950 4450
rect 3950 4398 4002 4450
rect 4002 4398 4004 4450
rect 3948 4396 4004 4398
rect 3836 4060 3892 4116
rect 3500 2940 3556 2996
rect 4620 6188 4676 6244
rect 4956 6076 5012 6132
rect 4844 5682 4900 5684
rect 4844 5630 4846 5682
rect 4846 5630 4898 5682
rect 4898 5630 4900 5682
rect 4844 5628 4900 5630
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4508 5292 4564 5348
rect 5292 6972 5348 7028
rect 5180 5740 5236 5796
rect 5292 6636 5348 6692
rect 5852 11900 5908 11956
rect 5740 10498 5796 10500
rect 5740 10446 5742 10498
rect 5742 10446 5794 10498
rect 5794 10446 5796 10498
rect 5740 10444 5796 10446
rect 5628 9996 5684 10052
rect 5628 8316 5684 8372
rect 5740 9324 5796 9380
rect 5628 8146 5684 8148
rect 5628 8094 5630 8146
rect 5630 8094 5682 8146
rect 5682 8094 5684 8146
rect 5628 8092 5684 8094
rect 6300 12124 6356 12180
rect 6076 11282 6132 11284
rect 6076 11230 6078 11282
rect 6078 11230 6130 11282
rect 6130 11230 6132 11282
rect 6076 11228 6132 11230
rect 6188 11170 6244 11172
rect 6188 11118 6190 11170
rect 6190 11118 6242 11170
rect 6242 11118 6244 11170
rect 6188 11116 6244 11118
rect 7196 11788 7252 11844
rect 6748 11116 6804 11172
rect 5964 9884 6020 9940
rect 6972 11004 7028 11060
rect 6076 9714 6132 9716
rect 6076 9662 6078 9714
rect 6078 9662 6130 9714
rect 6130 9662 6132 9714
rect 6076 9660 6132 9662
rect 6300 10722 6356 10724
rect 6300 10670 6302 10722
rect 6302 10670 6354 10722
rect 6354 10670 6356 10722
rect 6300 10668 6356 10670
rect 6860 10610 6916 10612
rect 6860 10558 6862 10610
rect 6862 10558 6914 10610
rect 6914 10558 6916 10610
rect 6860 10556 6916 10558
rect 6748 9996 6804 10052
rect 7644 11004 7700 11060
rect 7868 11004 7924 11060
rect 6076 9154 6132 9156
rect 6076 9102 6078 9154
rect 6078 9102 6130 9154
rect 6130 9102 6132 9154
rect 6076 9100 6132 9102
rect 5964 8540 6020 8596
rect 6300 9042 6356 9044
rect 6300 8990 6302 9042
rect 6302 8990 6354 9042
rect 6354 8990 6356 9042
rect 6300 8988 6356 8990
rect 7196 9436 7252 9492
rect 7084 9154 7140 9156
rect 7084 9102 7086 9154
rect 7086 9102 7138 9154
rect 7138 9102 7140 9154
rect 7084 9100 7140 9102
rect 6860 8876 6916 8932
rect 5852 8034 5908 8036
rect 5852 7982 5854 8034
rect 5854 7982 5906 8034
rect 5906 7982 5908 8034
rect 5852 7980 5908 7982
rect 5852 7250 5908 7252
rect 5852 7198 5854 7250
rect 5854 7198 5906 7250
rect 5906 7198 5908 7250
rect 5852 7196 5908 7198
rect 5740 7084 5796 7140
rect 6076 7084 6132 7140
rect 5628 6466 5684 6468
rect 5628 6414 5630 6466
rect 5630 6414 5682 6466
rect 5682 6414 5684 6466
rect 5628 6412 5684 6414
rect 5516 6018 5572 6020
rect 5516 5966 5518 6018
rect 5518 5966 5570 6018
rect 5570 5966 5572 6018
rect 5516 5964 5572 5966
rect 5964 6578 6020 6580
rect 5964 6526 5966 6578
rect 5966 6526 6018 6578
rect 6018 6526 6020 6578
rect 5964 6524 6020 6526
rect 5740 6018 5796 6020
rect 5740 5966 5742 6018
rect 5742 5966 5794 6018
rect 5794 5966 5796 6018
rect 5740 5964 5796 5966
rect 5292 5516 5348 5572
rect 5404 5180 5460 5236
rect 4620 5010 4676 5012
rect 4620 4958 4622 5010
rect 4622 4958 4674 5010
rect 4674 4958 4676 5010
rect 4620 4956 4676 4958
rect 5740 5122 5796 5124
rect 5740 5070 5742 5122
rect 5742 5070 5794 5122
rect 5794 5070 5796 5122
rect 5740 5068 5796 5070
rect 4956 4898 5012 4900
rect 4956 4846 4958 4898
rect 4958 4846 5010 4898
rect 5010 4846 5012 4898
rect 4956 4844 5012 4846
rect 4732 4562 4788 4564
rect 4732 4510 4734 4562
rect 4734 4510 4786 4562
rect 4786 4510 4788 4562
rect 4732 4508 4788 4510
rect 5852 4396 5908 4452
rect 5180 4172 5236 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4844 3500 4900 3556
rect 4172 3276 4228 3332
rect 7308 8988 7364 9044
rect 7420 9996 7476 10052
rect 8540 12684 8596 12740
rect 8092 11340 8148 11396
rect 8204 11788 8260 11844
rect 8428 11340 8484 11396
rect 7644 9548 7700 9604
rect 7420 8764 7476 8820
rect 6636 8034 6692 8036
rect 6636 7982 6638 8034
rect 6638 7982 6690 8034
rect 6690 7982 6692 8034
rect 6636 7980 6692 7982
rect 6748 7756 6804 7812
rect 7196 8092 7252 8148
rect 6972 7586 7028 7588
rect 6972 7534 6974 7586
rect 6974 7534 7026 7586
rect 7026 7534 7028 7586
rect 6972 7532 7028 7534
rect 7084 7980 7140 8036
rect 6524 7084 6580 7140
rect 6300 6972 6356 7028
rect 6524 6802 6580 6804
rect 6524 6750 6526 6802
rect 6526 6750 6578 6802
rect 6578 6750 6580 6802
rect 6524 6748 6580 6750
rect 6860 7362 6916 7364
rect 6860 7310 6862 7362
rect 6862 7310 6914 7362
rect 6914 7310 6916 7362
rect 6860 7308 6916 7310
rect 6636 6412 6692 6468
rect 6748 6130 6804 6132
rect 6748 6078 6750 6130
rect 6750 6078 6802 6130
rect 6802 6078 6804 6130
rect 6748 6076 6804 6078
rect 6972 6018 7028 6020
rect 6972 5966 6974 6018
rect 6974 5966 7026 6018
rect 7026 5966 7028 6018
rect 6972 5964 7028 5966
rect 6524 5906 6580 5908
rect 6524 5854 6526 5906
rect 6526 5854 6578 5906
rect 6578 5854 6580 5906
rect 6524 5852 6580 5854
rect 6300 5516 6356 5572
rect 7756 9042 7812 9044
rect 7756 8990 7758 9042
rect 7758 8990 7810 9042
rect 7810 8990 7812 9042
rect 7756 8988 7812 8990
rect 7980 9266 8036 9268
rect 7980 9214 7982 9266
rect 7982 9214 8034 9266
rect 8034 9214 8036 9266
rect 7980 9212 8036 9214
rect 7756 8540 7812 8596
rect 7868 8092 7924 8148
rect 7532 8034 7588 8036
rect 7532 7982 7534 8034
rect 7534 7982 7586 8034
rect 7586 7982 7588 8034
rect 7532 7980 7588 7982
rect 7420 7644 7476 7700
rect 7756 6636 7812 6692
rect 7308 5628 7364 5684
rect 6636 5180 6692 5236
rect 7868 5628 7924 5684
rect 7644 4956 7700 5012
rect 6860 4732 6916 4788
rect 7756 4844 7812 4900
rect 6076 4226 6132 4228
rect 6076 4174 6078 4226
rect 6078 4174 6130 4226
rect 6130 4174 6132 4226
rect 6076 4172 6132 4174
rect 7308 4226 7364 4228
rect 7308 4174 7310 4226
rect 7310 4174 7362 4226
rect 7362 4174 7364 4226
rect 7308 4172 7364 4174
rect 5964 4060 6020 4116
rect 8316 10610 8372 10612
rect 8316 10558 8318 10610
rect 8318 10558 8370 10610
rect 8370 10558 8372 10610
rect 8316 10556 8372 10558
rect 8988 13634 9044 13636
rect 8988 13582 8990 13634
rect 8990 13582 9042 13634
rect 9042 13582 9044 13634
rect 8988 13580 9044 13582
rect 8652 11788 8708 11844
rect 8652 11282 8708 11284
rect 8652 11230 8654 11282
rect 8654 11230 8706 11282
rect 8706 11230 8708 11282
rect 8652 11228 8708 11230
rect 8876 11004 8932 11060
rect 8988 10892 9044 10948
rect 8988 9884 9044 9940
rect 8764 9212 8820 9268
rect 9324 12236 9380 12292
rect 9436 12348 9492 12404
rect 9100 9212 9156 9268
rect 9212 9660 9268 9716
rect 8876 9154 8932 9156
rect 8876 9102 8878 9154
rect 8878 9102 8930 9154
rect 8930 9102 8932 9154
rect 8876 9100 8932 9102
rect 8092 8876 8148 8932
rect 8204 8316 8260 8372
rect 8652 8818 8708 8820
rect 8652 8766 8654 8818
rect 8654 8766 8706 8818
rect 8706 8766 8708 8818
rect 8652 8764 8708 8766
rect 8652 8428 8708 8484
rect 7980 5516 8036 5572
rect 8988 8930 9044 8932
rect 8988 8878 8990 8930
rect 8990 8878 9042 8930
rect 9042 8878 9044 8930
rect 8988 8876 9044 8878
rect 8876 8764 8932 8820
rect 9212 8764 9268 8820
rect 8876 7532 8932 7588
rect 9100 7868 9156 7924
rect 8652 7308 8708 7364
rect 8876 6412 8932 6468
rect 8428 5628 8484 5684
rect 8316 5516 8372 5572
rect 8988 5234 9044 5236
rect 8988 5182 8990 5234
rect 8990 5182 9042 5234
rect 9042 5182 9044 5234
rect 8988 5180 9044 5182
rect 9436 9884 9492 9940
rect 9436 8316 9492 8372
rect 9436 6748 9492 6804
rect 9324 6524 9380 6580
rect 11116 13804 11172 13860
rect 10332 13634 10388 13636
rect 10332 13582 10334 13634
rect 10334 13582 10386 13634
rect 10386 13582 10388 13634
rect 10332 13580 10388 13582
rect 9884 12460 9940 12516
rect 9884 12290 9940 12292
rect 9884 12238 9886 12290
rect 9886 12238 9938 12290
rect 9938 12238 9940 12290
rect 9884 12236 9940 12238
rect 9772 12012 9828 12068
rect 9660 11788 9716 11844
rect 10668 12738 10724 12740
rect 10668 12686 10670 12738
rect 10670 12686 10722 12738
rect 10722 12686 10724 12738
rect 10668 12684 10724 12686
rect 10220 12348 10276 12404
rect 10556 12124 10612 12180
rect 9884 11170 9940 11172
rect 9884 11118 9886 11170
rect 9886 11118 9938 11170
rect 9938 11118 9940 11170
rect 9884 11116 9940 11118
rect 10108 11452 10164 11508
rect 9884 10722 9940 10724
rect 9884 10670 9886 10722
rect 9886 10670 9938 10722
rect 9938 10670 9940 10722
rect 9884 10668 9940 10670
rect 10332 11116 10388 11172
rect 9996 10444 10052 10500
rect 9884 10386 9940 10388
rect 9884 10334 9886 10386
rect 9886 10334 9938 10386
rect 9938 10334 9940 10386
rect 9884 10332 9940 10334
rect 9772 9884 9828 9940
rect 9884 9266 9940 9268
rect 9884 9214 9886 9266
rect 9886 9214 9938 9266
rect 9938 9214 9940 9266
rect 9884 9212 9940 9214
rect 11116 12348 11172 12404
rect 11228 12796 11284 12852
rect 11004 12178 11060 12180
rect 11004 12126 11006 12178
rect 11006 12126 11058 12178
rect 11058 12126 11060 12178
rect 11004 12124 11060 12126
rect 10556 11676 10612 11732
rect 10108 9772 10164 9828
rect 10108 9154 10164 9156
rect 10108 9102 10110 9154
rect 10110 9102 10162 9154
rect 10162 9102 10164 9154
rect 10108 9100 10164 9102
rect 10220 8988 10276 9044
rect 9772 8652 9828 8708
rect 11116 11788 11172 11844
rect 10892 11228 10948 11284
rect 11004 11170 11060 11172
rect 11004 11118 11006 11170
rect 11006 11118 11058 11170
rect 11058 11118 11060 11170
rect 11004 11116 11060 11118
rect 18172 18508 18228 18564
rect 17276 17164 17332 17220
rect 15260 16882 15316 16884
rect 15260 16830 15262 16882
rect 15262 16830 15314 16882
rect 15314 16830 15316 16882
rect 15260 16828 15316 16830
rect 13356 15538 13412 15540
rect 13356 15486 13358 15538
rect 13358 15486 13410 15538
rect 13410 15486 13412 15538
rect 13356 15484 13412 15486
rect 14364 15484 14420 15540
rect 12572 15202 12628 15204
rect 12572 15150 12574 15202
rect 12574 15150 12626 15202
rect 12626 15150 12628 15202
rect 12572 15148 12628 15150
rect 13916 15202 13972 15204
rect 13916 15150 13918 15202
rect 13918 15150 13970 15202
rect 13970 15150 13972 15202
rect 13916 15148 13972 15150
rect 12012 13634 12068 13636
rect 12012 13582 12014 13634
rect 12014 13582 12066 13634
rect 12066 13582 12068 13634
rect 12012 13580 12068 13582
rect 11452 12738 11508 12740
rect 11452 12686 11454 12738
rect 11454 12686 11506 12738
rect 11506 12686 11508 12738
rect 11452 12684 11508 12686
rect 11452 11788 11508 11844
rect 11564 12460 11620 12516
rect 12012 12850 12068 12852
rect 12012 12798 12014 12850
rect 12014 12798 12066 12850
rect 12066 12798 12068 12850
rect 12012 12796 12068 12798
rect 12348 12572 12404 12628
rect 12908 13804 12964 13860
rect 12908 13634 12964 13636
rect 12908 13582 12910 13634
rect 12910 13582 12962 13634
rect 12962 13582 12964 13634
rect 12908 13580 12964 13582
rect 12796 12684 12852 12740
rect 12908 12572 12964 12628
rect 12460 12460 12516 12516
rect 11788 11676 11844 11732
rect 11676 11564 11732 11620
rect 12012 12124 12068 12180
rect 11676 11282 11732 11284
rect 11676 11230 11678 11282
rect 11678 11230 11730 11282
rect 11730 11230 11732 11282
rect 11676 11228 11732 11230
rect 11900 11170 11956 11172
rect 11900 11118 11902 11170
rect 11902 11118 11954 11170
rect 11954 11118 11956 11170
rect 11900 11116 11956 11118
rect 12572 12178 12628 12180
rect 12572 12126 12574 12178
rect 12574 12126 12626 12178
rect 12626 12126 12628 12178
rect 12572 12124 12628 12126
rect 12124 11340 12180 11396
rect 11564 9826 11620 9828
rect 11564 9774 11566 9826
rect 11566 9774 11618 9826
rect 11618 9774 11620 9826
rect 11564 9772 11620 9774
rect 10892 9660 10948 9716
rect 10556 8876 10612 8932
rect 9548 6412 9604 6468
rect 9660 8204 9716 8260
rect 9660 7308 9716 7364
rect 9660 6748 9716 6804
rect 10332 8428 10388 8484
rect 9996 7644 10052 7700
rect 10780 9212 10836 9268
rect 10668 8204 10724 8260
rect 10108 7586 10164 7588
rect 10108 7534 10110 7586
rect 10110 7534 10162 7586
rect 10162 7534 10164 7586
rect 10108 7532 10164 7534
rect 10668 7474 10724 7476
rect 10668 7422 10670 7474
rect 10670 7422 10722 7474
rect 10722 7422 10724 7474
rect 10668 7420 10724 7422
rect 9884 6636 9940 6692
rect 10444 6412 10500 6468
rect 10332 6188 10388 6244
rect 10220 5852 10276 5908
rect 9212 4620 9268 4676
rect 9100 4508 9156 4564
rect 10332 5740 10388 5796
rect 10556 5682 10612 5684
rect 10556 5630 10558 5682
rect 10558 5630 10610 5682
rect 10610 5630 10612 5682
rect 10556 5628 10612 5630
rect 10892 8316 10948 8372
rect 10780 4844 10836 4900
rect 10220 4732 10276 4788
rect 9772 3554 9828 3556
rect 9772 3502 9774 3554
rect 9774 3502 9826 3554
rect 9826 3502 9828 3554
rect 9772 3500 9828 3502
rect 11116 7196 11172 7252
rect 11564 8764 11620 8820
rect 11452 8316 11508 8372
rect 11900 9884 11956 9940
rect 12012 9100 12068 9156
rect 11676 8540 11732 8596
rect 11340 8204 11396 8260
rect 11564 6130 11620 6132
rect 11564 6078 11566 6130
rect 11566 6078 11618 6130
rect 11618 6078 11620 6130
rect 11564 6076 11620 6078
rect 11788 7362 11844 7364
rect 11788 7310 11790 7362
rect 11790 7310 11842 7362
rect 11842 7310 11844 7362
rect 11788 7308 11844 7310
rect 12124 8370 12180 8372
rect 12124 8318 12126 8370
rect 12126 8318 12178 8370
rect 12178 8318 12180 8370
rect 12124 8316 12180 8318
rect 12348 11788 12404 11844
rect 12460 11676 12516 11732
rect 12796 11676 12852 11732
rect 12460 10780 12516 10836
rect 12236 8204 12292 8260
rect 12908 11452 12964 11508
rect 13132 13804 13188 13860
rect 13356 13746 13412 13748
rect 13356 13694 13358 13746
rect 13358 13694 13410 13746
rect 13410 13694 13412 13746
rect 13356 13692 13412 13694
rect 13692 13692 13748 13748
rect 12908 10668 12964 10724
rect 12796 9714 12852 9716
rect 12796 9662 12798 9714
rect 12798 9662 12850 9714
rect 12850 9662 12852 9714
rect 12796 9660 12852 9662
rect 12572 9100 12628 9156
rect 12236 7644 12292 7700
rect 12460 8204 12516 8260
rect 12124 6076 12180 6132
rect 11340 5010 11396 5012
rect 11340 4958 11342 5010
rect 11342 4958 11394 5010
rect 11394 4958 11396 5010
rect 11340 4956 11396 4958
rect 11228 4732 11284 4788
rect 11116 4396 11172 4452
rect 12012 5010 12068 5012
rect 12012 4958 12014 5010
rect 12014 4958 12066 5010
rect 12066 4958 12068 5010
rect 12012 4956 12068 4958
rect 12572 5122 12628 5124
rect 12572 5070 12574 5122
rect 12574 5070 12626 5122
rect 12626 5070 12628 5122
rect 12572 5068 12628 5070
rect 12124 4898 12180 4900
rect 12124 4846 12126 4898
rect 12126 4846 12178 4898
rect 12178 4846 12180 4898
rect 12124 4844 12180 4846
rect 11900 4396 11956 4452
rect 12796 7308 12852 7364
rect 12796 6748 12852 6804
rect 13020 10780 13076 10836
rect 13468 12572 13524 12628
rect 13804 12738 13860 12740
rect 13804 12686 13806 12738
rect 13806 12686 13858 12738
rect 13858 12686 13860 12738
rect 13804 12684 13860 12686
rect 13580 12124 13636 12180
rect 13692 12572 13748 12628
rect 13132 9772 13188 9828
rect 13244 11340 13300 11396
rect 12684 4396 12740 4452
rect 13020 6636 13076 6692
rect 12908 5292 12964 5348
rect 13356 11228 13412 11284
rect 13356 5852 13412 5908
rect 13468 7644 13524 7700
rect 14252 13858 14308 13860
rect 14252 13806 14254 13858
rect 14254 13806 14306 13858
rect 14306 13806 14308 13858
rect 14252 13804 14308 13806
rect 13916 12572 13972 12628
rect 13692 11900 13748 11956
rect 13804 11676 13860 11732
rect 13916 11506 13972 11508
rect 13916 11454 13918 11506
rect 13918 11454 13970 11506
rect 13970 11454 13972 11506
rect 13916 11452 13972 11454
rect 13804 9884 13860 9940
rect 13916 11170 13972 11172
rect 13916 11118 13918 11170
rect 13918 11118 13970 11170
rect 13970 11118 13972 11170
rect 13916 11116 13972 11118
rect 13916 9660 13972 9716
rect 13580 5964 13636 6020
rect 13804 9548 13860 9604
rect 13468 5628 13524 5684
rect 13244 5068 13300 5124
rect 13692 5516 13748 5572
rect 13580 4396 13636 4452
rect 12908 4172 12964 4228
rect 13244 4060 13300 4116
rect 13244 3612 13300 3668
rect 14700 13692 14756 13748
rect 14588 13244 14644 13300
rect 14588 12908 14644 12964
rect 14364 12684 14420 12740
rect 14476 12572 14532 12628
rect 14252 12290 14308 12292
rect 14252 12238 14254 12290
rect 14254 12238 14306 12290
rect 14306 12238 14308 12290
rect 14252 12236 14308 12238
rect 14476 12124 14532 12180
rect 14476 11340 14532 11396
rect 14140 9660 14196 9716
rect 14028 8204 14084 8260
rect 14028 7084 14084 7140
rect 13916 6748 13972 6804
rect 13916 5628 13972 5684
rect 14028 4956 14084 5012
rect 14028 4508 14084 4564
rect 14476 11116 14532 11172
rect 14252 7644 14308 7700
rect 14252 6748 14308 6804
rect 14812 12572 14868 12628
rect 14924 13804 14980 13860
rect 14924 13580 14980 13636
rect 14700 11676 14756 11732
rect 14812 12348 14868 12404
rect 15260 14252 15316 14308
rect 15148 14140 15204 14196
rect 15148 13804 15204 13860
rect 15036 12908 15092 12964
rect 15148 12402 15204 12404
rect 15148 12350 15150 12402
rect 15150 12350 15202 12402
rect 15202 12350 15204 12402
rect 15148 12348 15204 12350
rect 14700 11282 14756 11284
rect 14700 11230 14702 11282
rect 14702 11230 14754 11282
rect 14754 11230 14756 11282
rect 14700 11228 14756 11230
rect 14812 8204 14868 8260
rect 14476 5906 14532 5908
rect 14476 5854 14478 5906
rect 14478 5854 14530 5906
rect 14530 5854 14532 5906
rect 14476 5852 14532 5854
rect 15708 15874 15764 15876
rect 15708 15822 15710 15874
rect 15710 15822 15762 15874
rect 15762 15822 15764 15874
rect 15708 15820 15764 15822
rect 15708 15484 15764 15540
rect 16044 15820 16100 15876
rect 15820 15202 15876 15204
rect 15820 15150 15822 15202
rect 15822 15150 15874 15202
rect 15874 15150 15876 15202
rect 15820 15148 15876 15150
rect 15484 14364 15540 14420
rect 15596 14306 15652 14308
rect 15596 14254 15598 14306
rect 15598 14254 15650 14306
rect 15650 14254 15652 14306
rect 15596 14252 15652 14254
rect 15708 13580 15764 13636
rect 16604 14812 16660 14868
rect 16492 14588 16548 14644
rect 16044 13634 16100 13636
rect 16044 13582 16046 13634
rect 16046 13582 16098 13634
rect 16098 13582 16100 13634
rect 16044 13580 16100 13582
rect 15484 12572 15540 12628
rect 15260 11788 15316 11844
rect 15372 11004 15428 11060
rect 15820 12402 15876 12404
rect 15820 12350 15822 12402
rect 15822 12350 15874 12402
rect 15874 12350 15876 12402
rect 15820 12348 15876 12350
rect 15820 12012 15876 12068
rect 15596 11900 15652 11956
rect 15820 11788 15876 11844
rect 15260 8428 15316 8484
rect 15148 8370 15204 8372
rect 15148 8318 15150 8370
rect 15150 8318 15202 8370
rect 15202 8318 15204 8370
rect 15148 8316 15204 8318
rect 15036 8258 15092 8260
rect 15036 8206 15038 8258
rect 15038 8206 15090 8258
rect 15090 8206 15092 8258
rect 15036 8204 15092 8206
rect 15372 6636 15428 6692
rect 15036 5906 15092 5908
rect 15036 5854 15038 5906
rect 15038 5854 15090 5906
rect 15090 5854 15092 5906
rect 15036 5852 15092 5854
rect 15596 11676 15652 11732
rect 15932 11564 15988 11620
rect 16044 11788 16100 11844
rect 15932 11394 15988 11396
rect 15932 11342 15934 11394
rect 15934 11342 15986 11394
rect 15986 11342 15988 11394
rect 15932 11340 15988 11342
rect 15596 8428 15652 8484
rect 15708 8316 15764 8372
rect 16044 7868 16100 7924
rect 16268 12738 16324 12740
rect 16268 12686 16270 12738
rect 16270 12686 16322 12738
rect 16322 12686 16324 12738
rect 16268 12684 16324 12686
rect 17052 14252 17108 14308
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 17948 15874 18004 15876
rect 17948 15822 17950 15874
rect 17950 15822 18002 15874
rect 18002 15822 18004 15874
rect 17948 15820 18004 15822
rect 18284 16882 18340 16884
rect 18284 16830 18286 16882
rect 18286 16830 18338 16882
rect 18338 16830 18340 16882
rect 18284 16828 18340 16830
rect 17500 15036 17556 15092
rect 17164 14140 17220 14196
rect 17388 14306 17444 14308
rect 17388 14254 17390 14306
rect 17390 14254 17442 14306
rect 17442 14254 17444 14306
rect 17388 14252 17444 14254
rect 16940 13970 16996 13972
rect 16940 13918 16942 13970
rect 16942 13918 16994 13970
rect 16994 13918 16996 13970
rect 16940 13916 16996 13918
rect 16828 12236 16884 12292
rect 17388 13692 17444 13748
rect 18172 14588 18228 14644
rect 17948 14476 18004 14532
rect 17948 13916 18004 13972
rect 17612 13580 17668 13636
rect 17276 12850 17332 12852
rect 17276 12798 17278 12850
rect 17278 12798 17330 12850
rect 17330 12798 17332 12850
rect 17276 12796 17332 12798
rect 16940 12124 16996 12180
rect 16716 11676 16772 11732
rect 16492 10668 16548 10724
rect 16604 11452 16660 11508
rect 16604 10556 16660 10612
rect 16604 10386 16660 10388
rect 16604 10334 16606 10386
rect 16606 10334 16658 10386
rect 16658 10334 16660 10386
rect 16604 10332 16660 10334
rect 17836 13692 17892 13748
rect 16940 11228 16996 11284
rect 16828 11116 16884 11172
rect 17276 11282 17332 11284
rect 17276 11230 17278 11282
rect 17278 11230 17330 11282
rect 17330 11230 17332 11282
rect 17276 11228 17332 11230
rect 17724 11788 17780 11844
rect 17500 10444 17556 10500
rect 17612 10668 17668 10724
rect 17948 10892 18004 10948
rect 17724 10220 17780 10276
rect 17724 9996 17780 10052
rect 17052 9100 17108 9156
rect 17500 9826 17556 9828
rect 17500 9774 17502 9826
rect 17502 9774 17554 9826
rect 17554 9774 17556 9826
rect 17500 9772 17556 9774
rect 17724 9660 17780 9716
rect 17276 8876 17332 8932
rect 17612 9324 17668 9380
rect 17388 8652 17444 8708
rect 16156 6748 16212 6804
rect 16604 6972 16660 7028
rect 17276 6914 17332 6916
rect 17276 6862 17278 6914
rect 17278 6862 17330 6914
rect 17330 6862 17332 6914
rect 17276 6860 17332 6862
rect 16716 6524 16772 6580
rect 16828 6636 16884 6692
rect 16828 6300 16884 6356
rect 17052 6636 17108 6692
rect 16828 6130 16884 6132
rect 16828 6078 16830 6130
rect 16830 6078 16882 6130
rect 16882 6078 16884 6130
rect 16828 6076 16884 6078
rect 16156 6018 16212 6020
rect 16156 5966 16158 6018
rect 16158 5966 16210 6018
rect 16210 5966 16212 6018
rect 16156 5964 16212 5966
rect 15820 5852 15876 5908
rect 15372 5628 15428 5684
rect 15036 5234 15092 5236
rect 15036 5182 15038 5234
rect 15038 5182 15090 5234
rect 15090 5182 15092 5234
rect 15036 5180 15092 5182
rect 15708 5180 15764 5236
rect 15596 4620 15652 4676
rect 14588 4172 14644 4228
rect 14252 3666 14308 3668
rect 14252 3614 14254 3666
rect 14254 3614 14306 3666
rect 14306 3614 14308 3666
rect 14252 3612 14308 3614
rect 14140 3500 14196 3556
rect 15484 4226 15540 4228
rect 15484 4174 15486 4226
rect 15486 4174 15538 4226
rect 15538 4174 15540 4226
rect 15484 4172 15540 4174
rect 16940 6018 16996 6020
rect 16940 5966 16942 6018
rect 16942 5966 16994 6018
rect 16994 5966 16996 6018
rect 16940 5964 16996 5966
rect 16828 5404 16884 5460
rect 17724 9266 17780 9268
rect 17724 9214 17726 9266
rect 17726 9214 17778 9266
rect 17778 9214 17780 9266
rect 17724 9212 17780 9214
rect 17948 8652 18004 8708
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 21980 39004 22036 39060
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 30044 27020 30100 27076
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 27020 24556 27076 24612
rect 25228 23884 25284 23940
rect 24780 23772 24836 23828
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 23324 22428 23380 22484
rect 18620 22092 18676 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21644 21868 21700 21924
rect 19628 21196 19684 21252
rect 19068 17948 19124 18004
rect 18732 17106 18788 17108
rect 18732 17054 18734 17106
rect 18734 17054 18786 17106
rect 18786 17054 18788 17106
rect 18732 17052 18788 17054
rect 18396 13468 18452 13524
rect 18508 16828 18564 16884
rect 19068 16770 19124 16772
rect 19068 16718 19070 16770
rect 19070 16718 19122 16770
rect 19122 16718 19124 16770
rect 19068 16716 19124 16718
rect 18732 16268 18788 16324
rect 18620 14924 18676 14980
rect 18620 13634 18676 13636
rect 18620 13582 18622 13634
rect 18622 13582 18674 13634
rect 18674 13582 18676 13634
rect 18620 13580 18676 13582
rect 18172 12124 18228 12180
rect 18284 12066 18340 12068
rect 18284 12014 18286 12066
rect 18286 12014 18338 12066
rect 18338 12014 18340 12066
rect 18284 12012 18340 12014
rect 18172 10722 18228 10724
rect 18172 10670 18174 10722
rect 18174 10670 18226 10722
rect 18226 10670 18228 10722
rect 18172 10668 18228 10670
rect 18284 10780 18340 10836
rect 18172 10332 18228 10388
rect 18396 9996 18452 10052
rect 18284 9436 18340 9492
rect 18396 9602 18452 9604
rect 18396 9550 18398 9602
rect 18398 9550 18450 9602
rect 18450 9550 18452 9602
rect 18396 9548 18452 9550
rect 18172 8930 18228 8932
rect 18172 8878 18174 8930
rect 18174 8878 18226 8930
rect 18226 8878 18228 8930
rect 18172 8876 18228 8878
rect 19180 16210 19236 16212
rect 19180 16158 19182 16210
rect 19182 16158 19234 16210
rect 19234 16158 19236 16210
rect 19180 16156 19236 16158
rect 18844 14252 18900 14308
rect 18732 12572 18788 12628
rect 18844 12684 18900 12740
rect 19068 14028 19124 14084
rect 19180 13692 19236 13748
rect 19516 17164 19572 17220
rect 19516 16940 19572 16996
rect 21084 20524 21140 20580
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20300 20188 20356 20244
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19852 18508 19908 18564
rect 20076 18338 20132 18340
rect 20076 18286 20078 18338
rect 20078 18286 20130 18338
rect 20130 18286 20132 18338
rect 20076 18284 20132 18286
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20188 17164 20244 17220
rect 20188 16604 20244 16660
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19964 15538 20020 15540
rect 19964 15486 19966 15538
rect 19966 15486 20018 15538
rect 20018 15486 20020 15538
rect 19964 15484 20020 15486
rect 19628 14476 19684 14532
rect 20076 14924 20132 14980
rect 19516 14364 19572 14420
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20188 14140 20244 14196
rect 19628 13916 19684 13972
rect 19404 13132 19460 13188
rect 19740 13692 19796 13748
rect 18844 12290 18900 12292
rect 18844 12238 18846 12290
rect 18846 12238 18898 12290
rect 18898 12238 18900 12290
rect 18844 12236 18900 12238
rect 18956 12124 19012 12180
rect 18732 10780 18788 10836
rect 18844 11340 18900 11396
rect 18732 10386 18788 10388
rect 18732 10334 18734 10386
rect 18734 10334 18786 10386
rect 18786 10334 18788 10386
rect 18732 10332 18788 10334
rect 18620 9602 18676 9604
rect 18620 9550 18622 9602
rect 18622 9550 18674 9602
rect 18674 9550 18676 9602
rect 18620 9548 18676 9550
rect 18508 9154 18564 9156
rect 18508 9102 18510 9154
rect 18510 9102 18562 9154
rect 18562 9102 18564 9154
rect 18508 9100 18564 9102
rect 18396 8428 18452 8484
rect 18060 8316 18116 8372
rect 18284 6972 18340 7028
rect 17612 5964 17668 6020
rect 17724 6524 17780 6580
rect 17164 4284 17220 4340
rect 17276 5180 17332 5236
rect 17836 6300 17892 6356
rect 18508 6636 18564 6692
rect 18620 7308 18676 7364
rect 18396 6466 18452 6468
rect 18396 6414 18398 6466
rect 18398 6414 18450 6466
rect 18450 6414 18452 6466
rect 18396 6412 18452 6414
rect 18284 6076 18340 6132
rect 17948 5906 18004 5908
rect 17948 5854 17950 5906
rect 17950 5854 18002 5906
rect 18002 5854 18004 5906
rect 17948 5852 18004 5854
rect 18508 5404 18564 5460
rect 18396 5234 18452 5236
rect 18396 5182 18398 5234
rect 18398 5182 18450 5234
rect 18450 5182 18452 5234
rect 18396 5180 18452 5182
rect 18844 9660 18900 9716
rect 19068 10722 19124 10724
rect 19068 10670 19070 10722
rect 19070 10670 19122 10722
rect 19122 10670 19124 10722
rect 19068 10668 19124 10670
rect 19180 9996 19236 10052
rect 19068 9826 19124 9828
rect 19068 9774 19070 9826
rect 19070 9774 19122 9826
rect 19122 9774 19124 9826
rect 19068 9772 19124 9774
rect 19180 9660 19236 9716
rect 18844 8876 18900 8932
rect 18956 9100 19012 9156
rect 19180 8930 19236 8932
rect 19180 8878 19182 8930
rect 19182 8878 19234 8930
rect 19234 8878 19236 8930
rect 19180 8876 19236 8878
rect 19180 8652 19236 8708
rect 19068 5964 19124 6020
rect 18732 4956 18788 5012
rect 18732 4396 18788 4452
rect 17836 3612 17892 3668
rect 17612 3554 17668 3556
rect 17612 3502 17614 3554
rect 17614 3502 17666 3554
rect 17666 3502 17668 3554
rect 17612 3500 17668 3502
rect 19404 12012 19460 12068
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19628 11900 19684 11956
rect 20188 11788 20244 11844
rect 19516 11452 19572 11508
rect 19964 11394 20020 11396
rect 19964 11342 19966 11394
rect 19966 11342 20018 11394
rect 20018 11342 20020 11394
rect 19964 11340 20020 11342
rect 19516 10892 19572 10948
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20076 10780 20132 10836
rect 19516 10668 19572 10724
rect 19964 10610 20020 10612
rect 19964 10558 19966 10610
rect 19966 10558 20018 10610
rect 20018 10558 20020 10610
rect 19964 10556 20020 10558
rect 19404 9938 19460 9940
rect 19404 9886 19406 9938
rect 19406 9886 19458 9938
rect 19458 9886 19460 9938
rect 19404 9884 19460 9886
rect 20188 10668 20244 10724
rect 19516 9436 19572 9492
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19516 8988 19572 9044
rect 19964 8258 20020 8260
rect 19964 8206 19966 8258
rect 19966 8206 20018 8258
rect 20018 8206 20020 8258
rect 19964 8204 20020 8206
rect 19740 8034 19796 8036
rect 19740 7982 19742 8034
rect 19742 7982 19794 8034
rect 19794 7982 19796 8034
rect 19740 7980 19796 7982
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20972 19740 21028 19796
rect 20748 19628 20804 19684
rect 20412 16322 20468 16324
rect 20412 16270 20414 16322
rect 20414 16270 20466 16322
rect 20466 16270 20468 16322
rect 20412 16268 20468 16270
rect 20860 18396 20916 18452
rect 20860 17778 20916 17780
rect 20860 17726 20862 17778
rect 20862 17726 20914 17778
rect 20914 17726 20916 17778
rect 20860 17724 20916 17726
rect 22988 21308 23044 21364
rect 22876 20748 22932 20804
rect 22876 20188 22932 20244
rect 26012 23548 26068 23604
rect 25564 22988 25620 23044
rect 26460 23100 26516 23156
rect 25564 22482 25620 22484
rect 25564 22430 25566 22482
rect 25566 22430 25618 22482
rect 25618 22430 25620 22482
rect 25564 22428 25620 22430
rect 24780 22092 24836 22148
rect 25564 22204 25620 22260
rect 24556 21474 24612 21476
rect 24556 21422 24558 21474
rect 24558 21422 24610 21474
rect 24610 21422 24612 21474
rect 24556 21420 24612 21422
rect 24108 21308 24164 21364
rect 23436 21084 23492 21140
rect 23884 20914 23940 20916
rect 23884 20862 23886 20914
rect 23886 20862 23938 20914
rect 23938 20862 23940 20914
rect 23884 20860 23940 20862
rect 24332 20690 24388 20692
rect 24332 20638 24334 20690
rect 24334 20638 24386 20690
rect 24386 20638 24388 20690
rect 24332 20636 24388 20638
rect 24668 20578 24724 20580
rect 24668 20526 24670 20578
rect 24670 20526 24722 20578
rect 24722 20526 24724 20578
rect 24668 20524 24724 20526
rect 25564 21474 25620 21476
rect 25564 21422 25566 21474
rect 25566 21422 25618 21474
rect 25618 21422 25620 21474
rect 25564 21420 25620 21422
rect 25788 20412 25844 20468
rect 22092 19906 22148 19908
rect 22092 19854 22094 19906
rect 22094 19854 22146 19906
rect 22146 19854 22148 19906
rect 22092 19852 22148 19854
rect 21644 18620 21700 18676
rect 21532 18396 21588 18452
rect 21308 18338 21364 18340
rect 21308 18286 21310 18338
rect 21310 18286 21362 18338
rect 21362 18286 21364 18338
rect 21308 18284 21364 18286
rect 21084 17164 21140 17220
rect 20860 16156 20916 16212
rect 20412 14028 20468 14084
rect 20860 14306 20916 14308
rect 20860 14254 20862 14306
rect 20862 14254 20914 14306
rect 20914 14254 20916 14306
rect 20860 14252 20916 14254
rect 20412 13692 20468 13748
rect 20412 12236 20468 12292
rect 20636 13244 20692 13300
rect 20524 11170 20580 11172
rect 20524 11118 20526 11170
rect 20526 11118 20578 11170
rect 20578 11118 20580 11170
rect 20524 11116 20580 11118
rect 20972 13692 21028 13748
rect 21308 17724 21364 17780
rect 21308 16940 21364 16996
rect 21756 18284 21812 18340
rect 22540 19516 22596 19572
rect 22540 19010 22596 19012
rect 22540 18958 22542 19010
rect 22542 18958 22594 19010
rect 22594 18958 22596 19010
rect 22540 18956 22596 18958
rect 22988 18732 23044 18788
rect 23660 19234 23716 19236
rect 23660 19182 23662 19234
rect 23662 19182 23714 19234
rect 23714 19182 23716 19234
rect 23660 19180 23716 19182
rect 23212 18508 23268 18564
rect 22092 17724 22148 17780
rect 21980 17164 22036 17220
rect 21756 16994 21812 16996
rect 21756 16942 21758 16994
rect 21758 16942 21810 16994
rect 21810 16942 21812 16994
rect 21756 16940 21812 16942
rect 23660 18508 23716 18564
rect 23772 17666 23828 17668
rect 23772 17614 23774 17666
rect 23774 17614 23826 17666
rect 23826 17614 23828 17666
rect 23772 17612 23828 17614
rect 22988 16940 23044 16996
rect 21644 15820 21700 15876
rect 21308 15426 21364 15428
rect 21308 15374 21310 15426
rect 21310 15374 21362 15426
rect 21362 15374 21364 15426
rect 21308 15372 21364 15374
rect 22428 16716 22484 16772
rect 22316 16156 22372 16212
rect 22204 15820 22260 15876
rect 21980 15372 22036 15428
rect 22652 16716 22708 16772
rect 22428 15372 22484 15428
rect 23324 16716 23380 16772
rect 24668 19906 24724 19908
rect 24668 19854 24670 19906
rect 24670 19854 24722 19906
rect 24722 19854 24724 19906
rect 24668 19852 24724 19854
rect 24220 19740 24276 19796
rect 24332 19068 24388 19124
rect 24108 18674 24164 18676
rect 24108 18622 24110 18674
rect 24110 18622 24162 18674
rect 24162 18622 24164 18674
rect 24108 18620 24164 18622
rect 24220 18396 24276 18452
rect 25004 19122 25060 19124
rect 25004 19070 25006 19122
rect 25006 19070 25058 19122
rect 25058 19070 25060 19122
rect 25004 19068 25060 19070
rect 24332 18562 24388 18564
rect 24332 18510 24334 18562
rect 24334 18510 24386 18562
rect 24386 18510 24388 18562
rect 24332 18508 24388 18510
rect 25228 19234 25284 19236
rect 25228 19182 25230 19234
rect 25230 19182 25282 19234
rect 25282 19182 25284 19234
rect 25228 19180 25284 19182
rect 25116 18956 25172 19012
rect 23996 17052 24052 17108
rect 24780 17612 24836 17668
rect 23212 16210 23268 16212
rect 23212 16158 23214 16210
rect 23214 16158 23266 16210
rect 23266 16158 23268 16210
rect 23212 16156 23268 16158
rect 23436 16044 23492 16100
rect 23100 15986 23156 15988
rect 23100 15934 23102 15986
rect 23102 15934 23154 15986
rect 23154 15934 23156 15986
rect 23100 15932 23156 15934
rect 23324 15372 23380 15428
rect 23436 15874 23492 15876
rect 23436 15822 23438 15874
rect 23438 15822 23490 15874
rect 23490 15822 23492 15874
rect 23436 15820 23492 15822
rect 24220 16268 24276 16324
rect 24668 16210 24724 16212
rect 24668 16158 24670 16210
rect 24670 16158 24722 16210
rect 24722 16158 24724 16210
rect 24668 16156 24724 16158
rect 24108 16098 24164 16100
rect 24108 16046 24110 16098
rect 24110 16046 24162 16098
rect 24162 16046 24164 16098
rect 24108 16044 24164 16046
rect 24332 16098 24388 16100
rect 24332 16046 24334 16098
rect 24334 16046 24386 16098
rect 24386 16046 24388 16098
rect 24332 16044 24388 16046
rect 24892 16604 24948 16660
rect 24780 16044 24836 16100
rect 24220 15820 24276 15876
rect 24668 15426 24724 15428
rect 24668 15374 24670 15426
rect 24670 15374 24722 15426
rect 24722 15374 24724 15426
rect 24668 15372 24724 15374
rect 25116 15372 25172 15428
rect 22988 15036 23044 15092
rect 23548 15036 23604 15092
rect 21420 14364 21476 14420
rect 21308 13858 21364 13860
rect 21308 13806 21310 13858
rect 21310 13806 21362 13858
rect 21362 13806 21364 13858
rect 21308 13804 21364 13806
rect 21084 13244 21140 13300
rect 20972 11788 21028 11844
rect 20524 8428 20580 8484
rect 19852 7644 19908 7700
rect 19852 6748 19908 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19852 6130 19908 6132
rect 19852 6078 19854 6130
rect 19854 6078 19906 6130
rect 19906 6078 19908 6130
rect 19852 6076 19908 6078
rect 19516 5068 19572 5124
rect 20524 7756 20580 7812
rect 20748 9884 20804 9940
rect 20860 9996 20916 10052
rect 20636 7532 20692 7588
rect 20636 7362 20692 7364
rect 20636 7310 20638 7362
rect 20638 7310 20690 7362
rect 20690 7310 20692 7362
rect 20636 7308 20692 7310
rect 20524 7084 20580 7140
rect 20748 6466 20804 6468
rect 20748 6414 20750 6466
rect 20750 6414 20802 6466
rect 20802 6414 20804 6466
rect 20748 6412 20804 6414
rect 20860 8316 20916 8372
rect 21756 14252 21812 14308
rect 21644 14028 21700 14084
rect 21532 13858 21588 13860
rect 21532 13806 21534 13858
rect 21534 13806 21586 13858
rect 21586 13806 21588 13858
rect 21532 13804 21588 13806
rect 21980 13020 22036 13076
rect 22316 13132 22372 13188
rect 21980 12850 22036 12852
rect 21980 12798 21982 12850
rect 21982 12798 22034 12850
rect 22034 12798 22036 12850
rect 21980 12796 22036 12798
rect 21756 11676 21812 11732
rect 22092 11564 22148 11620
rect 21196 8428 21252 8484
rect 21308 8092 21364 8148
rect 21644 10050 21700 10052
rect 21644 9998 21646 10050
rect 21646 9998 21698 10050
rect 21698 9998 21700 10050
rect 21644 9996 21700 9998
rect 21980 10108 22036 10164
rect 22204 11170 22260 11172
rect 22204 11118 22206 11170
rect 22206 11118 22258 11170
rect 22258 11118 22260 11170
rect 22204 11116 22260 11118
rect 22204 10780 22260 10836
rect 23212 13804 23268 13860
rect 22764 13580 22820 13636
rect 22652 13356 22708 13412
rect 22988 13074 23044 13076
rect 22988 13022 22990 13074
rect 22990 13022 23042 13074
rect 23042 13022 23044 13074
rect 22988 13020 23044 13022
rect 22652 12124 22708 12180
rect 22316 9996 22372 10052
rect 22092 9772 22148 9828
rect 22316 9826 22372 9828
rect 22316 9774 22318 9826
rect 22318 9774 22370 9826
rect 22370 9774 22372 9826
rect 22316 9772 22372 9774
rect 22540 9938 22596 9940
rect 22540 9886 22542 9938
rect 22542 9886 22594 9938
rect 22594 9886 22596 9938
rect 22540 9884 22596 9886
rect 22988 12796 23044 12852
rect 22876 11564 22932 11620
rect 22876 11004 22932 11060
rect 23436 13580 23492 13636
rect 25564 20130 25620 20132
rect 25564 20078 25566 20130
rect 25566 20078 25618 20130
rect 25618 20078 25620 20130
rect 25564 20076 25620 20078
rect 25564 17164 25620 17220
rect 26572 23042 26628 23044
rect 26572 22990 26574 23042
rect 26574 22990 26626 23042
rect 26626 22990 26628 23042
rect 26572 22988 26628 22990
rect 26236 21980 26292 22036
rect 26908 22146 26964 22148
rect 26908 22094 26910 22146
rect 26910 22094 26962 22146
rect 26962 22094 26964 22146
rect 26908 22092 26964 22094
rect 26908 21868 26964 21924
rect 26348 21532 26404 21588
rect 25900 19740 25956 19796
rect 26012 20018 26068 20020
rect 26012 19966 26014 20018
rect 26014 19966 26066 20018
rect 26066 19966 26068 20018
rect 26012 19964 26068 19966
rect 26236 20802 26292 20804
rect 26236 20750 26238 20802
rect 26238 20750 26290 20802
rect 26290 20750 26292 20802
rect 26236 20748 26292 20750
rect 26124 19852 26180 19908
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 25788 17890 25844 17892
rect 25788 17838 25790 17890
rect 25790 17838 25842 17890
rect 25842 17838 25844 17890
rect 25788 17836 25844 17838
rect 25452 16098 25508 16100
rect 25452 16046 25454 16098
rect 25454 16046 25506 16098
rect 25506 16046 25508 16098
rect 25452 16044 25508 16046
rect 25676 15372 25732 15428
rect 25228 15036 25284 15092
rect 25228 14364 25284 14420
rect 24220 14252 24276 14308
rect 23548 13356 23604 13412
rect 23660 13468 23716 13524
rect 23660 12178 23716 12180
rect 23660 12126 23662 12178
rect 23662 12126 23714 12178
rect 23714 12126 23716 12178
rect 23660 12124 23716 12126
rect 23212 11452 23268 11508
rect 22764 10220 22820 10276
rect 22428 9324 22484 9380
rect 22988 9436 23044 9492
rect 22316 9100 22372 9156
rect 21644 8876 21700 8932
rect 22428 8316 22484 8372
rect 22540 8988 22596 9044
rect 21420 7756 21476 7812
rect 21308 7308 21364 7364
rect 20300 5292 20356 5348
rect 19628 5010 19684 5012
rect 19628 4958 19630 5010
rect 19630 4958 19682 5010
rect 19682 4958 19684 5010
rect 19628 4956 19684 4958
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20860 5234 20916 5236
rect 20860 5182 20862 5234
rect 20862 5182 20914 5234
rect 20914 5182 20916 5234
rect 20860 5180 20916 5182
rect 21308 4226 21364 4228
rect 21308 4174 21310 4226
rect 21310 4174 21362 4226
rect 21362 4174 21364 4226
rect 21308 4172 21364 4174
rect 21420 6748 21476 6804
rect 21308 3948 21364 4004
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21532 6636 21588 6692
rect 21756 7868 21812 7924
rect 21532 5180 21588 5236
rect 21644 5068 21700 5124
rect 22092 7980 22148 8036
rect 21980 7756 22036 7812
rect 22988 9042 23044 9044
rect 22988 8990 22990 9042
rect 22990 8990 23042 9042
rect 23042 8990 23044 9042
rect 22988 8988 23044 8990
rect 23548 11788 23604 11844
rect 23884 11676 23940 11732
rect 23436 10722 23492 10724
rect 23436 10670 23438 10722
rect 23438 10670 23490 10722
rect 23490 10670 23492 10722
rect 23436 10668 23492 10670
rect 23212 9772 23268 9828
rect 23660 10332 23716 10388
rect 23100 8876 23156 8932
rect 22876 8316 22932 8372
rect 22204 6578 22260 6580
rect 22204 6526 22206 6578
rect 22206 6526 22258 6578
rect 22258 6526 22260 6578
rect 22204 6524 22260 6526
rect 22428 6412 22484 6468
rect 22764 6690 22820 6692
rect 22764 6638 22766 6690
rect 22766 6638 22818 6690
rect 22818 6638 22820 6690
rect 22764 6636 22820 6638
rect 22652 6076 22708 6132
rect 23100 7980 23156 8036
rect 23212 7084 23268 7140
rect 22988 6636 23044 6692
rect 23772 9826 23828 9828
rect 23772 9774 23774 9826
rect 23774 9774 23826 9826
rect 23826 9774 23828 9826
rect 23772 9772 23828 9774
rect 23548 9212 23604 9268
rect 23548 9042 23604 9044
rect 23548 8990 23550 9042
rect 23550 8990 23602 9042
rect 23602 8990 23604 9042
rect 23548 8988 23604 8990
rect 23660 8876 23716 8932
rect 23548 8428 23604 8484
rect 24444 13692 24500 13748
rect 24332 12684 24388 12740
rect 24332 11788 24388 11844
rect 23996 9714 24052 9716
rect 23996 9662 23998 9714
rect 23998 9662 24050 9714
rect 24050 9662 24052 9714
rect 23996 9660 24052 9662
rect 23996 9324 24052 9380
rect 23660 7474 23716 7476
rect 23660 7422 23662 7474
rect 23662 7422 23714 7474
rect 23714 7422 23716 7474
rect 23660 7420 23716 7422
rect 24108 9042 24164 9044
rect 24108 8990 24110 9042
rect 24110 8990 24162 9042
rect 24162 8990 24164 9042
rect 24108 8988 24164 8990
rect 24780 13692 24836 13748
rect 24556 13580 24612 13636
rect 24668 13356 24724 13412
rect 24668 10780 24724 10836
rect 24892 13356 24948 13412
rect 24892 12796 24948 12852
rect 24444 10332 24500 10388
rect 25004 10108 25060 10164
rect 24556 9324 24612 9380
rect 25452 13916 25508 13972
rect 25452 13692 25508 13748
rect 25340 12124 25396 12180
rect 24668 9100 24724 9156
rect 24780 9042 24836 9044
rect 24780 8990 24782 9042
rect 24782 8990 24834 9042
rect 24834 8990 24836 9042
rect 24780 8988 24836 8990
rect 24220 8764 24276 8820
rect 24668 8764 24724 8820
rect 24332 8652 24388 8708
rect 23100 6466 23156 6468
rect 23100 6414 23102 6466
rect 23102 6414 23154 6466
rect 23154 6414 23156 6466
rect 23100 6412 23156 6414
rect 23436 6412 23492 6468
rect 22988 6300 23044 6356
rect 22204 5740 22260 5796
rect 22204 4172 22260 4228
rect 23100 4844 23156 4900
rect 24108 6636 24164 6692
rect 23772 6188 23828 6244
rect 23660 5628 23716 5684
rect 23996 5964 24052 6020
rect 24668 8540 24724 8596
rect 24444 7362 24500 7364
rect 24444 7310 24446 7362
rect 24446 7310 24498 7362
rect 24498 7310 24500 7362
rect 24444 7308 24500 7310
rect 25228 8370 25284 8372
rect 25228 8318 25230 8370
rect 25230 8318 25282 8370
rect 25282 8318 25284 8370
rect 25228 8316 25284 8318
rect 25564 14812 25620 14868
rect 26124 18450 26180 18452
rect 26124 18398 26126 18450
rect 26126 18398 26178 18450
rect 26178 18398 26180 18450
rect 26124 18396 26180 18398
rect 26236 17836 26292 17892
rect 26012 17778 26068 17780
rect 26012 17726 26014 17778
rect 26014 17726 26066 17778
rect 26066 17726 26068 17778
rect 26012 17724 26068 17726
rect 26236 17388 26292 17444
rect 26684 21586 26740 21588
rect 26684 21534 26686 21586
rect 26686 21534 26738 21586
rect 26738 21534 26740 21586
rect 26684 21532 26740 21534
rect 26572 20690 26628 20692
rect 26572 20638 26574 20690
rect 26574 20638 26626 20690
rect 26626 20638 26628 20690
rect 26572 20636 26628 20638
rect 28028 24050 28084 24052
rect 28028 23998 28030 24050
rect 28030 23998 28082 24050
rect 28082 23998 28084 24050
rect 28028 23996 28084 23998
rect 36316 27020 36372 27076
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 33068 25228 33124 25284
rect 30492 24668 30548 24724
rect 28700 23212 28756 23268
rect 27804 22258 27860 22260
rect 27804 22206 27806 22258
rect 27806 22206 27858 22258
rect 27858 22206 27860 22258
rect 27804 22204 27860 22206
rect 27132 21644 27188 21700
rect 27020 20578 27076 20580
rect 27020 20526 27022 20578
rect 27022 20526 27074 20578
rect 27074 20526 27076 20578
rect 27020 20524 27076 20526
rect 27132 20076 27188 20132
rect 26908 19740 26964 19796
rect 27580 20524 27636 20580
rect 27356 19628 27412 19684
rect 27132 19404 27188 19460
rect 26572 18620 26628 18676
rect 27132 19010 27188 19012
rect 27132 18958 27134 19010
rect 27134 18958 27186 19010
rect 27186 18958 27188 19010
rect 27132 18956 27188 18958
rect 27132 18620 27188 18676
rect 26684 18396 26740 18452
rect 27020 18396 27076 18452
rect 26572 17554 26628 17556
rect 26572 17502 26574 17554
rect 26574 17502 26626 17554
rect 26626 17502 26628 17554
rect 26572 17500 26628 17502
rect 26684 17442 26740 17444
rect 26684 17390 26686 17442
rect 26686 17390 26738 17442
rect 26738 17390 26740 17442
rect 26684 17388 26740 17390
rect 26460 16940 26516 16996
rect 25900 16658 25956 16660
rect 25900 16606 25902 16658
rect 25902 16606 25954 16658
rect 25954 16606 25956 16658
rect 25900 16604 25956 16606
rect 25900 16098 25956 16100
rect 25900 16046 25902 16098
rect 25902 16046 25954 16098
rect 25954 16046 25956 16098
rect 25900 16044 25956 16046
rect 26348 16210 26404 16212
rect 26348 16158 26350 16210
rect 26350 16158 26402 16210
rect 26402 16158 26404 16210
rect 26348 16156 26404 16158
rect 26236 15708 26292 15764
rect 26012 15314 26068 15316
rect 26012 15262 26014 15314
rect 26014 15262 26066 15314
rect 26066 15262 26068 15314
rect 26012 15260 26068 15262
rect 26348 14812 26404 14868
rect 25900 14476 25956 14532
rect 26572 16828 26628 16884
rect 26572 14476 26628 14532
rect 25900 14306 25956 14308
rect 25900 14254 25902 14306
rect 25902 14254 25954 14306
rect 25954 14254 25956 14306
rect 25900 14252 25956 14254
rect 25676 13746 25732 13748
rect 25676 13694 25678 13746
rect 25678 13694 25730 13746
rect 25730 13694 25732 13746
rect 25676 13692 25732 13694
rect 25900 13746 25956 13748
rect 25900 13694 25902 13746
rect 25902 13694 25954 13746
rect 25954 13694 25956 13746
rect 25900 13692 25956 13694
rect 25788 13634 25844 13636
rect 25788 13582 25790 13634
rect 25790 13582 25842 13634
rect 25842 13582 25844 13634
rect 25788 13580 25844 13582
rect 26348 13746 26404 13748
rect 26348 13694 26350 13746
rect 26350 13694 26402 13746
rect 26402 13694 26404 13746
rect 26348 13692 26404 13694
rect 26236 13244 26292 13300
rect 26012 13020 26068 13076
rect 25900 12684 25956 12740
rect 25452 11452 25508 11508
rect 25452 10332 25508 10388
rect 25788 11340 25844 11396
rect 25900 11452 25956 11508
rect 25676 10444 25732 10500
rect 25564 10108 25620 10164
rect 25676 9996 25732 10052
rect 25564 9660 25620 9716
rect 25676 9324 25732 9380
rect 25676 8876 25732 8932
rect 24668 6748 24724 6804
rect 24780 7532 24836 7588
rect 24220 6188 24276 6244
rect 24220 5516 24276 5572
rect 23548 4956 23604 5012
rect 24220 5346 24276 5348
rect 24220 5294 24222 5346
rect 24222 5294 24274 5346
rect 24274 5294 24276 5346
rect 24220 5292 24276 5294
rect 23996 5180 24052 5236
rect 24220 4956 24276 5012
rect 24108 4844 24164 4900
rect 23996 4732 24052 4788
rect 22316 3948 22372 4004
rect 24108 4338 24164 4340
rect 24108 4286 24110 4338
rect 24110 4286 24162 4338
rect 24162 4286 24164 4338
rect 24108 4284 24164 4286
rect 23996 3724 24052 3780
rect 21532 3666 21588 3668
rect 21532 3614 21534 3666
rect 21534 3614 21586 3666
rect 21586 3614 21588 3666
rect 21532 3612 21588 3614
rect 22652 2940 22708 2996
rect 24220 3612 24276 3668
rect 24444 6076 24500 6132
rect 24444 5906 24500 5908
rect 24444 5854 24446 5906
rect 24446 5854 24498 5906
rect 24498 5854 24500 5906
rect 24444 5852 24500 5854
rect 24892 7308 24948 7364
rect 24892 6972 24948 7028
rect 24892 5852 24948 5908
rect 25004 6748 25060 6804
rect 25452 6690 25508 6692
rect 25452 6638 25454 6690
rect 25454 6638 25506 6690
rect 25506 6638 25508 6690
rect 25452 6636 25508 6638
rect 25900 10722 25956 10724
rect 25900 10670 25902 10722
rect 25902 10670 25954 10722
rect 25954 10670 25956 10722
rect 25900 10668 25956 10670
rect 26124 10780 26180 10836
rect 25900 10444 25956 10500
rect 26012 10332 26068 10388
rect 25788 8652 25844 8708
rect 26124 9154 26180 9156
rect 26124 9102 26126 9154
rect 26126 9102 26178 9154
rect 26178 9102 26180 9154
rect 26124 9100 26180 9102
rect 26124 8204 26180 8260
rect 26572 12796 26628 12852
rect 26908 17554 26964 17556
rect 26908 17502 26910 17554
rect 26910 17502 26962 17554
rect 26962 17502 26964 17554
rect 26908 17500 26964 17502
rect 27020 16882 27076 16884
rect 27020 16830 27022 16882
rect 27022 16830 27074 16882
rect 27074 16830 27076 16882
rect 27020 16828 27076 16830
rect 27356 17890 27412 17892
rect 27356 17838 27358 17890
rect 27358 17838 27410 17890
rect 27410 17838 27412 17890
rect 27356 17836 27412 17838
rect 27468 17554 27524 17556
rect 27468 17502 27470 17554
rect 27470 17502 27522 17554
rect 27522 17502 27524 17554
rect 27468 17500 27524 17502
rect 27244 17276 27300 17332
rect 27244 16940 27300 16996
rect 27468 16492 27524 16548
rect 27356 16380 27412 16436
rect 27020 15708 27076 15764
rect 26908 15596 26964 15652
rect 27132 15538 27188 15540
rect 27132 15486 27134 15538
rect 27134 15486 27186 15538
rect 27186 15486 27188 15538
rect 27132 15484 27188 15486
rect 26796 15314 26852 15316
rect 26796 15262 26798 15314
rect 26798 15262 26850 15314
rect 26850 15262 26852 15314
rect 26796 15260 26852 15262
rect 27244 15148 27300 15204
rect 27356 15932 27412 15988
rect 27020 15036 27076 15092
rect 27468 15314 27524 15316
rect 27468 15262 27470 15314
rect 27470 15262 27522 15314
rect 27522 15262 27524 15314
rect 27468 15260 27524 15262
rect 27132 14530 27188 14532
rect 27132 14478 27134 14530
rect 27134 14478 27186 14530
rect 27186 14478 27188 14530
rect 27132 14476 27188 14478
rect 27244 14306 27300 14308
rect 27244 14254 27246 14306
rect 27246 14254 27298 14306
rect 27298 14254 27300 14306
rect 27244 14252 27300 14254
rect 27244 13916 27300 13972
rect 26908 13746 26964 13748
rect 26908 13694 26910 13746
rect 26910 13694 26962 13746
rect 26962 13694 26964 13746
rect 26908 13692 26964 13694
rect 26796 13020 26852 13076
rect 27132 13074 27188 13076
rect 27132 13022 27134 13074
rect 27134 13022 27186 13074
rect 27186 13022 27188 13074
rect 27132 13020 27188 13022
rect 26684 12572 26740 12628
rect 27356 13746 27412 13748
rect 27356 13694 27358 13746
rect 27358 13694 27410 13746
rect 27410 13694 27412 13746
rect 27356 13692 27412 13694
rect 28028 21474 28084 21476
rect 28028 21422 28030 21474
rect 28030 21422 28082 21474
rect 28082 21422 28084 21474
rect 28028 21420 28084 21422
rect 27804 20972 27860 21028
rect 27916 20412 27972 20468
rect 27804 20018 27860 20020
rect 27804 19966 27806 20018
rect 27806 19966 27858 20018
rect 27858 19966 27860 20018
rect 27804 19964 27860 19966
rect 27692 19628 27748 19684
rect 28588 22876 28644 22932
rect 28140 20972 28196 21028
rect 28252 22540 28308 22596
rect 28812 22428 28868 22484
rect 28364 20300 28420 20356
rect 28028 19404 28084 19460
rect 28140 19964 28196 20020
rect 28140 19292 28196 19348
rect 28252 19628 28308 19684
rect 28028 19180 28084 19236
rect 28140 18508 28196 18564
rect 28028 17388 28084 17444
rect 27804 16380 27860 16436
rect 29484 22482 29540 22484
rect 29484 22430 29486 22482
rect 29486 22430 29538 22482
rect 29538 22430 29540 22482
rect 29484 22428 29540 22430
rect 29372 21868 29428 21924
rect 28812 21810 28868 21812
rect 28812 21758 28814 21810
rect 28814 21758 28866 21810
rect 28866 21758 28868 21810
rect 28812 21756 28868 21758
rect 28700 20690 28756 20692
rect 28700 20638 28702 20690
rect 28702 20638 28754 20690
rect 28754 20638 28756 20690
rect 28700 20636 28756 20638
rect 28588 20524 28644 20580
rect 29708 23154 29764 23156
rect 29708 23102 29710 23154
rect 29710 23102 29762 23154
rect 29762 23102 29764 23154
rect 29708 23100 29764 23102
rect 30044 22876 30100 22932
rect 29596 20860 29652 20916
rect 29932 22652 29988 22708
rect 30044 22316 30100 22372
rect 30604 24610 30660 24612
rect 30604 24558 30606 24610
rect 30606 24558 30658 24610
rect 30658 24558 30660 24610
rect 30604 24556 30660 24558
rect 30492 23548 30548 23604
rect 30828 23100 30884 23156
rect 30492 22540 30548 22596
rect 30716 22540 30772 22596
rect 30492 22370 30548 22372
rect 30492 22318 30494 22370
rect 30494 22318 30546 22370
rect 30546 22318 30548 22370
rect 30492 22316 30548 22318
rect 30268 22204 30324 22260
rect 30604 22204 30660 22260
rect 29484 20578 29540 20580
rect 29484 20526 29486 20578
rect 29486 20526 29538 20578
rect 29538 20526 29540 20578
rect 29484 20524 29540 20526
rect 28588 19628 28644 19684
rect 29148 19628 29204 19684
rect 28588 18508 28644 18564
rect 29148 19292 29204 19348
rect 28476 16940 28532 16996
rect 28588 18060 28644 18116
rect 28924 18060 28980 18116
rect 28364 16828 28420 16884
rect 28476 16716 28532 16772
rect 28252 16380 28308 16436
rect 28364 16492 28420 16548
rect 28140 15484 28196 15540
rect 28252 16098 28308 16100
rect 28252 16046 28254 16098
rect 28254 16046 28306 16098
rect 28306 16046 28308 16098
rect 28252 16044 28308 16046
rect 28028 15036 28084 15092
rect 28364 15932 28420 15988
rect 28028 14252 28084 14308
rect 28028 13580 28084 13636
rect 27356 13020 27412 13076
rect 26348 10108 26404 10164
rect 27132 11954 27188 11956
rect 27132 11902 27134 11954
rect 27134 11902 27186 11954
rect 27186 11902 27188 11954
rect 27132 11900 27188 11902
rect 26908 11676 26964 11732
rect 26684 11564 26740 11620
rect 26572 10722 26628 10724
rect 26572 10670 26574 10722
rect 26574 10670 26626 10722
rect 26626 10670 26628 10722
rect 26572 10668 26628 10670
rect 26684 9996 26740 10052
rect 26796 10220 26852 10276
rect 26684 9324 26740 9380
rect 28924 16716 28980 16772
rect 28588 16044 28644 16100
rect 28476 15708 28532 15764
rect 28588 15372 28644 15428
rect 28476 15036 28532 15092
rect 28476 14812 28532 14868
rect 28812 15202 28868 15204
rect 28812 15150 28814 15202
rect 28814 15150 28866 15202
rect 28866 15150 28868 15202
rect 28812 15148 28868 15150
rect 28700 14700 28756 14756
rect 28588 14476 28644 14532
rect 28812 14418 28868 14420
rect 28812 14366 28814 14418
rect 28814 14366 28866 14418
rect 28866 14366 28868 14418
rect 28812 14364 28868 14366
rect 28588 14028 28644 14084
rect 28476 13858 28532 13860
rect 28476 13806 28478 13858
rect 28478 13806 28530 13858
rect 28530 13806 28532 13858
rect 28476 13804 28532 13806
rect 28364 13356 28420 13412
rect 28588 13356 28644 13412
rect 28252 13244 28308 13300
rect 27692 12850 27748 12852
rect 27692 12798 27694 12850
rect 27694 12798 27746 12850
rect 27746 12798 27748 12850
rect 27692 12796 27748 12798
rect 27468 11676 27524 11732
rect 27580 12290 27636 12292
rect 27580 12238 27582 12290
rect 27582 12238 27634 12290
rect 27634 12238 27636 12290
rect 27580 12236 27636 12238
rect 27244 11228 27300 11284
rect 27580 11004 27636 11060
rect 27356 9826 27412 9828
rect 27356 9774 27358 9826
rect 27358 9774 27410 9826
rect 27410 9774 27412 9826
rect 27356 9772 27412 9774
rect 27468 9714 27524 9716
rect 27468 9662 27470 9714
rect 27470 9662 27522 9714
rect 27522 9662 27524 9714
rect 27468 9660 27524 9662
rect 27916 11900 27972 11956
rect 27916 11228 27972 11284
rect 27916 10780 27972 10836
rect 28140 12738 28196 12740
rect 28140 12686 28142 12738
rect 28142 12686 28194 12738
rect 28194 12686 28196 12738
rect 28140 12684 28196 12686
rect 28476 13132 28532 13188
rect 28364 12850 28420 12852
rect 28364 12798 28366 12850
rect 28366 12798 28418 12850
rect 28418 12798 28420 12850
rect 28364 12796 28420 12798
rect 28252 12290 28308 12292
rect 28252 12238 28254 12290
rect 28254 12238 28306 12290
rect 28306 12238 28308 12290
rect 28252 12236 28308 12238
rect 28252 11954 28308 11956
rect 28252 11902 28254 11954
rect 28254 11902 28306 11954
rect 28306 11902 28308 11954
rect 28252 11900 28308 11902
rect 28476 11900 28532 11956
rect 28700 12908 28756 12964
rect 29372 18956 29428 19012
rect 29260 18172 29316 18228
rect 29036 14588 29092 14644
rect 28924 14252 28980 14308
rect 29148 14476 29204 14532
rect 30156 19906 30212 19908
rect 30156 19854 30158 19906
rect 30158 19854 30210 19906
rect 30210 19854 30212 19906
rect 30156 19852 30212 19854
rect 30716 20300 30772 20356
rect 30604 20188 30660 20244
rect 30044 19740 30100 19796
rect 29932 19292 29988 19348
rect 29596 19180 29652 19236
rect 29932 19010 29988 19012
rect 29932 18958 29934 19010
rect 29934 18958 29986 19010
rect 29986 18958 29988 19010
rect 29932 18956 29988 18958
rect 31388 22652 31444 22708
rect 31724 23212 31780 23268
rect 31500 22540 31556 22596
rect 30940 21868 30996 21924
rect 31276 22092 31332 22148
rect 31612 21756 31668 21812
rect 31836 23100 31892 23156
rect 35756 24668 35812 24724
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35756 24050 35812 24052
rect 35756 23998 35758 24050
rect 35758 23998 35810 24050
rect 35810 23998 35812 24050
rect 35756 23996 35812 23998
rect 34188 23938 34244 23940
rect 34188 23886 34190 23938
rect 34190 23886 34242 23938
rect 34242 23886 34244 23938
rect 35980 24556 36036 24612
rect 34188 23884 34244 23886
rect 31276 21644 31332 21700
rect 30828 19740 30884 19796
rect 30716 18844 30772 18900
rect 29484 18396 29540 18452
rect 29372 18060 29428 18116
rect 29596 16492 29652 16548
rect 29708 18396 29764 18452
rect 29484 15596 29540 15652
rect 29596 15484 29652 15540
rect 31724 21644 31780 21700
rect 31836 22204 31892 22260
rect 31724 21474 31780 21476
rect 31724 21422 31726 21474
rect 31726 21422 31778 21474
rect 31778 21422 31780 21474
rect 31724 21420 31780 21422
rect 31836 20578 31892 20580
rect 31836 20526 31838 20578
rect 31838 20526 31890 20578
rect 31890 20526 31892 20578
rect 31836 20524 31892 20526
rect 31836 20242 31892 20244
rect 31836 20190 31838 20242
rect 31838 20190 31890 20242
rect 31890 20190 31892 20242
rect 31836 20188 31892 20190
rect 31052 19906 31108 19908
rect 31052 19854 31054 19906
rect 31054 19854 31106 19906
rect 31106 19854 31108 19906
rect 31052 19852 31108 19854
rect 31052 18956 31108 19012
rect 30940 18508 30996 18564
rect 29820 17164 29876 17220
rect 30044 18060 30100 18116
rect 30268 17666 30324 17668
rect 30268 17614 30270 17666
rect 30270 17614 30322 17666
rect 30322 17614 30324 17666
rect 30268 17612 30324 17614
rect 30156 17442 30212 17444
rect 30156 17390 30158 17442
rect 30158 17390 30210 17442
rect 30210 17390 30212 17442
rect 30156 17388 30212 17390
rect 30604 18338 30660 18340
rect 30604 18286 30606 18338
rect 30606 18286 30658 18338
rect 30658 18286 30660 18338
rect 30604 18284 30660 18286
rect 31052 18338 31108 18340
rect 31052 18286 31054 18338
rect 31054 18286 31106 18338
rect 31106 18286 31108 18338
rect 31052 18284 31108 18286
rect 30492 18226 30548 18228
rect 30492 18174 30494 18226
rect 30494 18174 30546 18226
rect 30546 18174 30548 18226
rect 30492 18172 30548 18174
rect 30380 16940 30436 16996
rect 29932 16770 29988 16772
rect 29932 16718 29934 16770
rect 29934 16718 29986 16770
rect 29986 16718 29988 16770
rect 29932 16716 29988 16718
rect 29820 15874 29876 15876
rect 29820 15822 29822 15874
rect 29822 15822 29874 15874
rect 29874 15822 29876 15874
rect 29820 15820 29876 15822
rect 29484 15426 29540 15428
rect 29484 15374 29486 15426
rect 29486 15374 29538 15426
rect 29538 15374 29540 15426
rect 29484 15372 29540 15374
rect 29372 15314 29428 15316
rect 29372 15262 29374 15314
rect 29374 15262 29426 15314
rect 29426 15262 29428 15314
rect 29372 15260 29428 15262
rect 29708 15314 29764 15316
rect 29708 15262 29710 15314
rect 29710 15262 29762 15314
rect 29762 15262 29764 15314
rect 29708 15260 29764 15262
rect 29484 15148 29540 15204
rect 29036 14140 29092 14196
rect 28364 10892 28420 10948
rect 27804 10108 27860 10164
rect 28028 10556 28084 10612
rect 27692 9938 27748 9940
rect 27692 9886 27694 9938
rect 27694 9886 27746 9938
rect 27746 9886 27748 9938
rect 27692 9884 27748 9886
rect 27132 9324 27188 9380
rect 27244 9266 27300 9268
rect 27244 9214 27246 9266
rect 27246 9214 27298 9266
rect 27298 9214 27300 9266
rect 27244 9212 27300 9214
rect 26236 8764 26292 8820
rect 26796 8540 26852 8596
rect 26460 7980 26516 8036
rect 25788 7420 25844 7476
rect 25228 6578 25284 6580
rect 25228 6526 25230 6578
rect 25230 6526 25282 6578
rect 25282 6526 25284 6578
rect 25228 6524 25284 6526
rect 26908 7756 26964 7812
rect 25564 6466 25620 6468
rect 25564 6414 25566 6466
rect 25566 6414 25618 6466
rect 25618 6414 25620 6466
rect 25564 6412 25620 6414
rect 25564 6130 25620 6132
rect 25564 6078 25566 6130
rect 25566 6078 25618 6130
rect 25618 6078 25620 6130
rect 25564 6076 25620 6078
rect 25228 5068 25284 5124
rect 25340 5628 25396 5684
rect 24780 4956 24836 5012
rect 24892 4508 24948 4564
rect 24892 4172 24948 4228
rect 24668 2828 24724 2884
rect 25564 5234 25620 5236
rect 25564 5182 25566 5234
rect 25566 5182 25618 5234
rect 25618 5182 25620 5234
rect 25564 5180 25620 5182
rect 25452 4396 25508 4452
rect 25004 3388 25060 3444
rect 25004 3276 25060 3332
rect 26348 6300 26404 6356
rect 25788 5852 25844 5908
rect 26348 5906 26404 5908
rect 26348 5854 26350 5906
rect 26350 5854 26402 5906
rect 26402 5854 26404 5906
rect 26348 5852 26404 5854
rect 27020 6690 27076 6692
rect 27020 6638 27022 6690
rect 27022 6638 27074 6690
rect 27074 6638 27076 6690
rect 27020 6636 27076 6638
rect 27132 6524 27188 6580
rect 26684 5852 26740 5908
rect 26124 5740 26180 5796
rect 26572 5516 26628 5572
rect 26796 5404 26852 5460
rect 26124 5292 26180 5348
rect 26012 4562 26068 4564
rect 26012 4510 26014 4562
rect 26014 4510 26066 4562
rect 26066 4510 26068 4562
rect 26012 4508 26068 4510
rect 26572 4396 26628 4452
rect 27020 5516 27076 5572
rect 26908 4956 26964 5012
rect 26460 4338 26516 4340
rect 26460 4286 26462 4338
rect 26462 4286 26514 4338
rect 26514 4286 26516 4338
rect 26460 4284 26516 4286
rect 26348 3724 26404 3780
rect 24892 2716 24948 2772
rect 25788 3388 25844 3444
rect 26908 3500 26964 3556
rect 27468 7756 27524 7812
rect 27356 5964 27412 6020
rect 27132 5180 27188 5236
rect 27804 9154 27860 9156
rect 27804 9102 27806 9154
rect 27806 9102 27858 9154
rect 27858 9102 27860 9154
rect 27804 9100 27860 9102
rect 27916 9042 27972 9044
rect 27916 8990 27918 9042
rect 27918 8990 27970 9042
rect 27970 8990 27972 9042
rect 27916 8988 27972 8990
rect 28364 10722 28420 10724
rect 28364 10670 28366 10722
rect 28366 10670 28418 10722
rect 28418 10670 28420 10722
rect 28364 10668 28420 10670
rect 28140 9772 28196 9828
rect 28252 8876 28308 8932
rect 28700 11506 28756 11508
rect 28700 11454 28702 11506
rect 28702 11454 28754 11506
rect 28754 11454 28756 11506
rect 28700 11452 28756 11454
rect 28924 11452 28980 11508
rect 28700 11004 28756 11060
rect 28700 10332 28756 10388
rect 28588 9602 28644 9604
rect 28588 9550 28590 9602
rect 28590 9550 28642 9602
rect 28642 9550 28644 9602
rect 28588 9548 28644 9550
rect 28476 9212 28532 9268
rect 28588 9154 28644 9156
rect 28588 9102 28590 9154
rect 28590 9102 28642 9154
rect 28642 9102 28644 9154
rect 28588 9100 28644 9102
rect 28364 8540 28420 8596
rect 28812 9660 28868 9716
rect 28924 9996 28980 10052
rect 28700 7868 28756 7924
rect 27916 7586 27972 7588
rect 27916 7534 27918 7586
rect 27918 7534 27970 7586
rect 27970 7534 27972 7586
rect 27916 7532 27972 7534
rect 27692 7308 27748 7364
rect 27916 7084 27972 7140
rect 28140 7420 28196 7476
rect 27916 6466 27972 6468
rect 27916 6414 27918 6466
rect 27918 6414 27970 6466
rect 27970 6414 27972 6466
rect 27916 6412 27972 6414
rect 27580 5906 27636 5908
rect 27580 5854 27582 5906
rect 27582 5854 27634 5906
rect 27634 5854 27636 5906
rect 27580 5852 27636 5854
rect 27468 5404 27524 5460
rect 27468 5068 27524 5124
rect 27804 5516 27860 5572
rect 28476 7474 28532 7476
rect 28476 7422 28478 7474
rect 28478 7422 28530 7474
rect 28530 7422 28532 7474
rect 28476 7420 28532 7422
rect 28588 7362 28644 7364
rect 28588 7310 28590 7362
rect 28590 7310 28642 7362
rect 28642 7310 28644 7362
rect 28588 7308 28644 7310
rect 28812 7308 28868 7364
rect 28812 7084 28868 7140
rect 28364 5852 28420 5908
rect 28476 5964 28532 6020
rect 28252 5794 28308 5796
rect 28252 5742 28254 5794
rect 28254 5742 28306 5794
rect 28306 5742 28308 5794
rect 28252 5740 28308 5742
rect 28364 5346 28420 5348
rect 28364 5294 28366 5346
rect 28366 5294 28418 5346
rect 28418 5294 28420 5346
rect 28364 5292 28420 5294
rect 27580 3554 27636 3556
rect 27580 3502 27582 3554
rect 27582 3502 27634 3554
rect 27634 3502 27636 3554
rect 27580 3500 27636 3502
rect 28140 4508 28196 4564
rect 26684 3388 26740 3444
rect 28588 5404 28644 5460
rect 28812 5180 28868 5236
rect 29708 14476 29764 14532
rect 29596 14028 29652 14084
rect 29260 13468 29316 13524
rect 29372 13580 29428 13636
rect 29148 12178 29204 12180
rect 29148 12126 29150 12178
rect 29150 12126 29202 12178
rect 29202 12126 29204 12178
rect 29148 12124 29204 12126
rect 29148 10780 29204 10836
rect 30044 16492 30100 16548
rect 30492 17948 30548 18004
rect 31164 18060 31220 18116
rect 30940 17778 30996 17780
rect 30940 17726 30942 17778
rect 30942 17726 30994 17778
rect 30994 17726 30996 17778
rect 30940 17724 30996 17726
rect 31388 19740 31444 19796
rect 32508 23548 32564 23604
rect 33292 23714 33348 23716
rect 33292 23662 33294 23714
rect 33294 23662 33346 23714
rect 33346 23662 33348 23714
rect 33292 23660 33348 23662
rect 32172 23212 32228 23268
rect 32508 23266 32564 23268
rect 32508 23214 32510 23266
rect 32510 23214 32562 23266
rect 32562 23214 32564 23266
rect 32508 23212 32564 23214
rect 33404 23212 33460 23268
rect 32620 22988 32676 23044
rect 32508 22316 32564 22372
rect 33516 23042 33572 23044
rect 33516 22990 33518 23042
rect 33518 22990 33570 23042
rect 33570 22990 33572 23042
rect 33516 22988 33572 22990
rect 35308 23714 35364 23716
rect 35308 23662 35310 23714
rect 35310 23662 35362 23714
rect 35362 23662 35364 23714
rect 35308 23660 35364 23662
rect 35084 23100 35140 23156
rect 33852 22988 33908 23044
rect 33964 22876 34020 22932
rect 34188 22988 34244 23044
rect 32172 21810 32228 21812
rect 32172 21758 32174 21810
rect 32174 21758 32226 21810
rect 32226 21758 32228 21810
rect 32172 21756 32228 21758
rect 32060 19852 32116 19908
rect 31948 19628 32004 19684
rect 31276 17724 31332 17780
rect 31500 18956 31556 19012
rect 31612 18844 31668 18900
rect 32284 19404 32340 19460
rect 31948 18732 32004 18788
rect 32284 19180 32340 19236
rect 31948 18060 32004 18116
rect 31500 17612 31556 17668
rect 31612 17948 31668 18004
rect 31052 17554 31108 17556
rect 31052 17502 31054 17554
rect 31054 17502 31106 17554
rect 31106 17502 31108 17554
rect 31052 17500 31108 17502
rect 30604 17164 30660 17220
rect 31276 17442 31332 17444
rect 31276 17390 31278 17442
rect 31278 17390 31330 17442
rect 31330 17390 31332 17442
rect 31276 17388 31332 17390
rect 31500 17388 31556 17444
rect 30716 16492 30772 16548
rect 31388 16994 31444 16996
rect 31388 16942 31390 16994
rect 31390 16942 31442 16994
rect 31442 16942 31444 16994
rect 31388 16940 31444 16942
rect 30940 16044 30996 16100
rect 31276 16604 31332 16660
rect 31724 17164 31780 17220
rect 32060 17164 32116 17220
rect 31724 16604 31780 16660
rect 31500 15986 31556 15988
rect 31500 15934 31502 15986
rect 31502 15934 31554 15986
rect 31554 15934 31556 15986
rect 31500 15932 31556 15934
rect 30044 15820 30100 15876
rect 30156 15708 30212 15764
rect 29932 13804 29988 13860
rect 29820 13468 29876 13524
rect 30380 15538 30436 15540
rect 30380 15486 30382 15538
rect 30382 15486 30434 15538
rect 30434 15486 30436 15538
rect 30380 15484 30436 15486
rect 30268 15260 30324 15316
rect 30604 15538 30660 15540
rect 30604 15486 30606 15538
rect 30606 15486 30658 15538
rect 30658 15486 30660 15538
rect 30604 15484 30660 15486
rect 31388 15484 31444 15540
rect 30716 15314 30772 15316
rect 30716 15262 30718 15314
rect 30718 15262 30770 15314
rect 30770 15262 30772 15314
rect 30716 15260 30772 15262
rect 31500 15148 31556 15204
rect 30492 14476 30548 14532
rect 30828 14812 30884 14868
rect 30604 14418 30660 14420
rect 30604 14366 30606 14418
rect 30606 14366 30658 14418
rect 30658 14366 30660 14418
rect 30604 14364 30660 14366
rect 30492 14306 30548 14308
rect 30492 14254 30494 14306
rect 30494 14254 30546 14306
rect 30546 14254 30548 14306
rect 30492 14252 30548 14254
rect 30492 13804 30548 13860
rect 30156 12962 30212 12964
rect 30156 12910 30158 12962
rect 30158 12910 30210 12962
rect 30210 12910 30212 12962
rect 30156 12908 30212 12910
rect 30380 12908 30436 12964
rect 29596 12178 29652 12180
rect 29596 12126 29598 12178
rect 29598 12126 29650 12178
rect 29650 12126 29652 12178
rect 29596 12124 29652 12126
rect 29932 12572 29988 12628
rect 29820 12348 29876 12404
rect 29708 11676 29764 11732
rect 29036 8540 29092 8596
rect 29036 6076 29092 6132
rect 29820 11116 29876 11172
rect 29596 9996 29652 10052
rect 29372 9772 29428 9828
rect 29260 9212 29316 9268
rect 29596 9772 29652 9828
rect 29708 10892 29764 10948
rect 29596 9212 29652 9268
rect 29820 10108 29876 10164
rect 29596 8876 29652 8932
rect 29484 8540 29540 8596
rect 30380 12124 30436 12180
rect 30604 12796 30660 12852
rect 31276 14754 31332 14756
rect 31276 14702 31278 14754
rect 31278 14702 31330 14754
rect 31330 14702 31332 14754
rect 31276 14700 31332 14702
rect 31836 16380 31892 16436
rect 31836 16098 31892 16100
rect 31836 16046 31838 16098
rect 31838 16046 31890 16098
rect 31890 16046 31892 16098
rect 31836 16044 31892 16046
rect 32172 17106 32228 17108
rect 32172 17054 32174 17106
rect 32174 17054 32226 17106
rect 32226 17054 32228 17106
rect 32172 17052 32228 17054
rect 32396 18396 32452 18452
rect 32620 21308 32676 21364
rect 32620 20524 32676 20580
rect 32620 20188 32676 20244
rect 33740 22146 33796 22148
rect 33740 22094 33742 22146
rect 33742 22094 33794 22146
rect 33794 22094 33796 22146
rect 33740 22092 33796 22094
rect 32844 20188 32900 20244
rect 34300 21980 34356 22036
rect 33740 21756 33796 21812
rect 33516 20914 33572 20916
rect 33516 20862 33518 20914
rect 33518 20862 33570 20914
rect 33570 20862 33572 20914
rect 33516 20860 33572 20862
rect 33068 19964 33124 20020
rect 32620 19740 32676 19796
rect 32620 18620 32676 18676
rect 32508 17666 32564 17668
rect 32508 17614 32510 17666
rect 32510 17614 32562 17666
rect 32562 17614 32564 17666
rect 32508 17612 32564 17614
rect 33516 20018 33572 20020
rect 33516 19966 33518 20018
rect 33518 19966 33570 20018
rect 33570 19966 33572 20018
rect 33516 19964 33572 19966
rect 33628 19852 33684 19908
rect 34524 21980 34580 22036
rect 34300 21756 34356 21812
rect 34076 21586 34132 21588
rect 34076 21534 34078 21586
rect 34078 21534 34130 21586
rect 34130 21534 34132 21586
rect 34076 21532 34132 21534
rect 34300 20860 34356 20916
rect 33964 20578 34020 20580
rect 33964 20526 33966 20578
rect 33966 20526 34018 20578
rect 34018 20526 34020 20578
rect 33964 20524 34020 20526
rect 34300 20524 34356 20580
rect 34412 20018 34468 20020
rect 34412 19966 34414 20018
rect 34414 19966 34466 20018
rect 34466 19966 34468 20018
rect 34412 19964 34468 19966
rect 33964 19906 34020 19908
rect 33964 19854 33966 19906
rect 33966 19854 34018 19906
rect 34018 19854 34020 19906
rect 33964 19852 34020 19854
rect 33740 19404 33796 19460
rect 33516 19180 33572 19236
rect 32732 18284 32788 18340
rect 32844 19010 32900 19012
rect 32844 18958 32846 19010
rect 32846 18958 32898 19010
rect 32898 18958 32900 19010
rect 32844 18956 32900 18958
rect 32620 17164 32676 17220
rect 32396 16994 32452 16996
rect 32396 16942 32398 16994
rect 32398 16942 32450 16994
rect 32450 16942 32452 16994
rect 32396 16940 32452 16942
rect 32508 16044 32564 16100
rect 32732 16828 32788 16884
rect 32284 15596 32340 15652
rect 32620 15596 32676 15652
rect 32172 15372 32228 15428
rect 32284 15314 32340 15316
rect 32284 15262 32286 15314
rect 32286 15262 32338 15314
rect 32338 15262 32340 15314
rect 32284 15260 32340 15262
rect 32508 15260 32564 15316
rect 32396 15148 32452 15204
rect 31052 13020 31108 13076
rect 30716 12684 30772 12740
rect 30716 12460 30772 12516
rect 31612 12850 31668 12852
rect 31612 12798 31614 12850
rect 31614 12798 31666 12850
rect 31666 12798 31668 12850
rect 31612 12796 31668 12798
rect 31500 12684 31556 12740
rect 30940 12460 30996 12516
rect 31612 12348 31668 12404
rect 30940 12178 30996 12180
rect 30940 12126 30942 12178
rect 30942 12126 30994 12178
rect 30994 12126 30996 12178
rect 30940 12124 30996 12126
rect 30828 12012 30884 12068
rect 30044 11676 30100 11732
rect 30604 11732 30660 11788
rect 30044 11004 30100 11060
rect 31052 12012 31108 12068
rect 31500 12012 31556 12068
rect 31164 11954 31220 11956
rect 31164 11902 31166 11954
rect 31166 11902 31218 11954
rect 31218 11902 31220 11954
rect 31164 11900 31220 11902
rect 30828 11170 30884 11172
rect 30828 11118 30830 11170
rect 30830 11118 30882 11170
rect 30882 11118 30884 11170
rect 30828 11116 30884 11118
rect 30268 10050 30324 10052
rect 30268 9998 30270 10050
rect 30270 9998 30322 10050
rect 30322 9998 30324 10050
rect 30268 9996 30324 9998
rect 30044 9938 30100 9940
rect 30044 9886 30046 9938
rect 30046 9886 30098 9938
rect 30098 9886 30100 9938
rect 30044 9884 30100 9886
rect 30156 9548 30212 9604
rect 29596 8370 29652 8372
rect 29596 8318 29598 8370
rect 29598 8318 29650 8370
rect 29650 8318 29652 8370
rect 29596 8316 29652 8318
rect 29260 7084 29316 7140
rect 29372 7644 29428 7700
rect 29260 6018 29316 6020
rect 29260 5966 29262 6018
rect 29262 5966 29314 6018
rect 29314 5966 29316 6018
rect 29260 5964 29316 5966
rect 29148 5292 29204 5348
rect 29708 7980 29764 8036
rect 29708 7698 29764 7700
rect 29708 7646 29710 7698
rect 29710 7646 29762 7698
rect 29762 7646 29764 7698
rect 29708 7644 29764 7646
rect 29596 7420 29652 7476
rect 29820 6860 29876 6916
rect 29932 6972 29988 7028
rect 29932 6748 29988 6804
rect 30604 9938 30660 9940
rect 30604 9886 30606 9938
rect 30606 9886 30658 9938
rect 30658 9886 30660 9938
rect 30604 9884 30660 9886
rect 30828 9660 30884 9716
rect 30492 8370 30548 8372
rect 30492 8318 30494 8370
rect 30494 8318 30546 8370
rect 30546 8318 30548 8370
rect 30492 8316 30548 8318
rect 30604 8034 30660 8036
rect 30604 7982 30606 8034
rect 30606 7982 30658 8034
rect 30658 7982 30660 8034
rect 30604 7980 30660 7982
rect 31164 11732 31220 11788
rect 31164 11340 31220 11396
rect 31388 10892 31444 10948
rect 31388 10722 31444 10724
rect 31388 10670 31390 10722
rect 31390 10670 31442 10722
rect 31442 10670 31444 10722
rect 31388 10668 31444 10670
rect 31500 10610 31556 10612
rect 31500 10558 31502 10610
rect 31502 10558 31554 10610
rect 31554 10558 31556 10610
rect 31500 10556 31556 10558
rect 31388 10220 31444 10276
rect 31164 9884 31220 9940
rect 31052 9602 31108 9604
rect 31052 9550 31054 9602
rect 31054 9550 31106 9602
rect 31106 9550 31108 9602
rect 31052 9548 31108 9550
rect 31276 9548 31332 9604
rect 30940 7868 30996 7924
rect 31164 8988 31220 9044
rect 30492 7644 30548 7700
rect 30604 7756 30660 7812
rect 30492 7474 30548 7476
rect 30492 7422 30494 7474
rect 30494 7422 30546 7474
rect 30546 7422 30548 7474
rect 30492 7420 30548 7422
rect 30828 7474 30884 7476
rect 30828 7422 30830 7474
rect 30830 7422 30882 7474
rect 30882 7422 30884 7474
rect 30828 7420 30884 7422
rect 30604 7308 30660 7364
rect 31388 9042 31444 9044
rect 31388 8990 31390 9042
rect 31390 8990 31442 9042
rect 31442 8990 31444 9042
rect 31388 8988 31444 8990
rect 31612 9826 31668 9828
rect 31612 9774 31614 9826
rect 31614 9774 31666 9826
rect 31666 9774 31668 9826
rect 31612 9772 31668 9774
rect 32172 14924 32228 14980
rect 32060 14364 32116 14420
rect 32844 16604 32900 16660
rect 32956 18338 33012 18340
rect 32956 18286 32958 18338
rect 32958 18286 33010 18338
rect 33010 18286 33012 18338
rect 32956 18284 33012 18286
rect 32844 16098 32900 16100
rect 32844 16046 32846 16098
rect 32846 16046 32898 16098
rect 32898 16046 32900 16098
rect 32844 16044 32900 16046
rect 34188 19234 34244 19236
rect 34188 19182 34190 19234
rect 34190 19182 34242 19234
rect 34242 19182 34244 19234
rect 34188 19180 34244 19182
rect 33292 19010 33348 19012
rect 33292 18958 33294 19010
rect 33294 18958 33346 19010
rect 33346 18958 33348 19010
rect 33292 18956 33348 18958
rect 33068 17388 33124 17444
rect 34076 18338 34132 18340
rect 34076 18286 34078 18338
rect 34078 18286 34130 18338
rect 34130 18286 34132 18338
rect 34076 18284 34132 18286
rect 33628 17612 33684 17668
rect 34076 18060 34132 18116
rect 33740 16940 33796 16996
rect 33292 16492 33348 16548
rect 33404 16156 33460 16212
rect 33628 16156 33684 16212
rect 32956 15932 33012 15988
rect 32844 15596 32900 15652
rect 32620 14530 32676 14532
rect 32620 14478 32622 14530
rect 32622 14478 32674 14530
rect 32674 14478 32676 14530
rect 32620 14476 32676 14478
rect 32172 14028 32228 14084
rect 32060 13634 32116 13636
rect 32060 13582 32062 13634
rect 32062 13582 32114 13634
rect 32114 13582 32116 13634
rect 32060 13580 32116 13582
rect 31948 12572 32004 12628
rect 32060 13020 32116 13076
rect 31836 10892 31892 10948
rect 32844 13916 32900 13972
rect 32508 13858 32564 13860
rect 32508 13806 32510 13858
rect 32510 13806 32562 13858
rect 32562 13806 32564 13858
rect 32508 13804 32564 13806
rect 32732 13692 32788 13748
rect 32396 13468 32452 13524
rect 33068 13356 33124 13412
rect 32956 11676 33012 11732
rect 33068 12236 33124 12292
rect 31948 9548 32004 9604
rect 32060 9436 32116 9492
rect 31388 8370 31444 8372
rect 31388 8318 31390 8370
rect 31390 8318 31442 8370
rect 31442 8318 31444 8370
rect 31388 8316 31444 8318
rect 31724 8540 31780 8596
rect 32732 11452 32788 11508
rect 32284 11004 32340 11060
rect 32844 11394 32900 11396
rect 32844 11342 32846 11394
rect 32846 11342 32898 11394
rect 32898 11342 32900 11394
rect 32844 11340 32900 11342
rect 33516 15314 33572 15316
rect 33516 15262 33518 15314
rect 33518 15262 33570 15314
rect 33570 15262 33572 15314
rect 33516 15260 33572 15262
rect 33852 16380 33908 16436
rect 33740 15260 33796 15316
rect 33516 14700 33572 14756
rect 33292 14588 33348 14644
rect 33628 14588 33684 14644
rect 33180 11340 33236 11396
rect 33292 13692 33348 13748
rect 32620 10834 32676 10836
rect 32620 10782 32622 10834
rect 32622 10782 32674 10834
rect 32674 10782 32676 10834
rect 32620 10780 32676 10782
rect 32508 10444 32564 10500
rect 32732 10332 32788 10388
rect 32172 9212 32228 9268
rect 32284 9042 32340 9044
rect 32284 8990 32286 9042
rect 32286 8990 32338 9042
rect 32338 8990 32340 9042
rect 32284 8988 32340 8990
rect 32060 8428 32116 8484
rect 31276 7756 31332 7812
rect 33628 14028 33684 14084
rect 33516 13020 33572 13076
rect 33628 13580 33684 13636
rect 34076 15260 34132 15316
rect 33964 15148 34020 15204
rect 34524 19180 34580 19236
rect 34524 18844 34580 18900
rect 34412 16882 34468 16884
rect 34412 16830 34414 16882
rect 34414 16830 34466 16882
rect 34466 16830 34468 16882
rect 34412 16828 34468 16830
rect 34636 17276 34692 17332
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22316 35140 22372
rect 35532 22146 35588 22148
rect 35532 22094 35534 22146
rect 35534 22094 35586 22146
rect 35586 22094 35588 22146
rect 35532 22092 35588 22094
rect 35084 21980 35140 22036
rect 34860 20300 34916 20356
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35868 21980 35924 22036
rect 35756 21868 35812 21924
rect 35756 20914 35812 20916
rect 35756 20862 35758 20914
rect 35758 20862 35810 20914
rect 35810 20862 35812 20914
rect 35756 20860 35812 20862
rect 35532 20524 35588 20580
rect 35868 20524 35924 20580
rect 34972 19964 35028 20020
rect 35084 19852 35140 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 18338 34916 18340
rect 34860 18286 34862 18338
rect 34862 18286 34914 18338
rect 34914 18286 34916 18338
rect 34860 18284 34916 18286
rect 34972 18226 35028 18228
rect 34972 18174 34974 18226
rect 34974 18174 35026 18226
rect 35026 18174 35028 18226
rect 34972 18172 35028 18174
rect 34748 17164 34804 17220
rect 34972 16156 35028 16212
rect 34412 15874 34468 15876
rect 34412 15822 34414 15874
rect 34414 15822 34466 15874
rect 34466 15822 34468 15874
rect 34412 15820 34468 15822
rect 34300 14418 34356 14420
rect 34300 14366 34302 14418
rect 34302 14366 34354 14418
rect 34354 14366 34356 14418
rect 34300 14364 34356 14366
rect 33852 13970 33908 13972
rect 33852 13918 33854 13970
rect 33854 13918 33906 13970
rect 33906 13918 33908 13970
rect 33852 13916 33908 13918
rect 33964 13356 34020 13412
rect 33852 13244 33908 13300
rect 33852 12178 33908 12180
rect 33852 12126 33854 12178
rect 33854 12126 33906 12178
rect 33906 12126 33908 12178
rect 33852 12124 33908 12126
rect 33964 13020 34020 13076
rect 33740 11564 33796 11620
rect 33292 10332 33348 10388
rect 33516 11228 33572 11284
rect 33740 10722 33796 10724
rect 33740 10670 33742 10722
rect 33742 10670 33794 10722
rect 33794 10670 33796 10722
rect 33740 10668 33796 10670
rect 33628 10610 33684 10612
rect 33628 10558 33630 10610
rect 33630 10558 33682 10610
rect 33682 10558 33684 10610
rect 33628 10556 33684 10558
rect 34300 13746 34356 13748
rect 34300 13694 34302 13746
rect 34302 13694 34354 13746
rect 34354 13694 34356 13746
rect 34300 13692 34356 13694
rect 34748 15986 34804 15988
rect 34748 15934 34750 15986
rect 34750 15934 34802 15986
rect 34802 15934 34804 15986
rect 34748 15932 34804 15934
rect 34524 14364 34580 14420
rect 34636 15484 34692 15540
rect 34860 15260 34916 15316
rect 34860 14812 34916 14868
rect 35756 19516 35812 19572
rect 35532 19180 35588 19236
rect 35420 18338 35476 18340
rect 35420 18286 35422 18338
rect 35422 18286 35474 18338
rect 35474 18286 35476 18338
rect 35420 18284 35476 18286
rect 35756 19010 35812 19012
rect 35756 18958 35758 19010
rect 35758 18958 35810 19010
rect 35810 18958 35812 19010
rect 35756 18956 35812 18958
rect 35644 18732 35700 18788
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35308 16156 35364 16212
rect 35868 18508 35924 18564
rect 43260 25228 43316 25284
rect 38444 24780 38500 24836
rect 36876 24050 36932 24052
rect 36876 23998 36878 24050
rect 36878 23998 36930 24050
rect 36930 23998 36932 24050
rect 36876 23996 36932 23998
rect 37548 23996 37604 24052
rect 36428 22652 36484 22708
rect 36540 22540 36596 22596
rect 36092 20860 36148 20916
rect 36204 20412 36260 20468
rect 36316 20300 36372 20356
rect 36204 19740 36260 19796
rect 35980 18172 36036 18228
rect 35420 15986 35476 15988
rect 35420 15934 35422 15986
rect 35422 15934 35474 15986
rect 35474 15934 35476 15986
rect 35420 15932 35476 15934
rect 35644 16380 35700 16436
rect 35644 15708 35700 15764
rect 35756 16156 35812 16212
rect 35644 15538 35700 15540
rect 35644 15486 35646 15538
rect 35646 15486 35698 15538
rect 35698 15486 35700 15538
rect 35644 15484 35700 15486
rect 35532 15314 35588 15316
rect 35532 15262 35534 15314
rect 35534 15262 35586 15314
rect 35586 15262 35588 15314
rect 35532 15260 35588 15262
rect 35644 15148 35700 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34972 14140 35028 14196
rect 34748 13580 34804 13636
rect 34188 11900 34244 11956
rect 34300 12290 34356 12292
rect 34300 12238 34302 12290
rect 34302 12238 34354 12290
rect 34354 12238 34356 12290
rect 34300 12236 34356 12238
rect 34188 11282 34244 11284
rect 34188 11230 34190 11282
rect 34190 11230 34242 11282
rect 34242 11230 34244 11282
rect 34188 11228 34244 11230
rect 34524 12290 34580 12292
rect 34524 12238 34526 12290
rect 34526 12238 34578 12290
rect 34578 12238 34580 12290
rect 34524 12236 34580 12238
rect 34412 11788 34468 11844
rect 34412 11452 34468 11508
rect 34524 11676 34580 11732
rect 34076 10892 34132 10948
rect 34300 10834 34356 10836
rect 34300 10782 34302 10834
rect 34302 10782 34354 10834
rect 34354 10782 34356 10834
rect 34300 10780 34356 10782
rect 34636 10892 34692 10948
rect 34524 10556 34580 10612
rect 33516 9436 33572 9492
rect 34300 10108 34356 10164
rect 33740 9324 33796 9380
rect 33964 9996 34020 10052
rect 33852 9266 33908 9268
rect 33852 9214 33854 9266
rect 33854 9214 33906 9266
rect 33906 9214 33908 9266
rect 33852 9212 33908 9214
rect 33628 8540 33684 8596
rect 33404 8370 33460 8372
rect 33404 8318 33406 8370
rect 33406 8318 33458 8370
rect 33458 8318 33460 8370
rect 33404 8316 33460 8318
rect 31612 7868 31668 7924
rect 32508 7756 32564 7812
rect 29708 6578 29764 6580
rect 29708 6526 29710 6578
rect 29710 6526 29762 6578
rect 29762 6526 29764 6578
rect 29708 6524 29764 6526
rect 29932 6300 29988 6356
rect 29372 5628 29428 5684
rect 29036 4620 29092 4676
rect 29260 3666 29316 3668
rect 29260 3614 29262 3666
rect 29262 3614 29314 3666
rect 29314 3614 29316 3666
rect 29260 3612 29316 3614
rect 30940 6578 30996 6580
rect 30940 6526 30942 6578
rect 30942 6526 30994 6578
rect 30994 6526 30996 6578
rect 30940 6524 30996 6526
rect 31276 6578 31332 6580
rect 31276 6526 31278 6578
rect 31278 6526 31330 6578
rect 31330 6526 31332 6578
rect 31276 6524 31332 6526
rect 30940 5906 30996 5908
rect 30940 5854 30942 5906
rect 30942 5854 30994 5906
rect 30994 5854 30996 5906
rect 30940 5852 30996 5854
rect 31052 5794 31108 5796
rect 31052 5742 31054 5794
rect 31054 5742 31106 5794
rect 31106 5742 31108 5794
rect 31052 5740 31108 5742
rect 30492 5516 30548 5572
rect 31052 5234 31108 5236
rect 31052 5182 31054 5234
rect 31054 5182 31106 5234
rect 31106 5182 31108 5234
rect 31052 5180 31108 5182
rect 30828 4956 30884 5012
rect 30044 4396 30100 4452
rect 30716 4450 30772 4452
rect 30716 4398 30718 4450
rect 30718 4398 30770 4450
rect 30770 4398 30772 4450
rect 30716 4396 30772 4398
rect 29932 4338 29988 4340
rect 29932 4286 29934 4338
rect 29934 4286 29986 4338
rect 29986 4286 29988 4338
rect 29932 4284 29988 4286
rect 25788 1596 25844 1652
rect 30268 3442 30324 3444
rect 30268 3390 30270 3442
rect 30270 3390 30322 3442
rect 30322 3390 30324 3442
rect 30268 3388 30324 3390
rect 29372 2604 29428 2660
rect 31500 5906 31556 5908
rect 31500 5854 31502 5906
rect 31502 5854 31554 5906
rect 31554 5854 31556 5906
rect 31500 5852 31556 5854
rect 31276 5404 31332 5460
rect 31388 5516 31444 5572
rect 31724 5740 31780 5796
rect 31836 5628 31892 5684
rect 32284 7250 32340 7252
rect 32284 7198 32286 7250
rect 32286 7198 32338 7250
rect 32338 7198 32340 7250
rect 32284 7196 32340 7198
rect 32060 5740 32116 5796
rect 33740 7980 33796 8036
rect 33068 7868 33124 7924
rect 32060 5404 32116 5460
rect 31836 4172 31892 4228
rect 32172 5180 32228 5236
rect 32732 6130 32788 6132
rect 32732 6078 32734 6130
rect 32734 6078 32786 6130
rect 32786 6078 32788 6130
rect 32732 6076 32788 6078
rect 32396 5906 32452 5908
rect 32396 5854 32398 5906
rect 32398 5854 32450 5906
rect 32450 5854 32452 5906
rect 32396 5852 32452 5854
rect 32620 5682 32676 5684
rect 32620 5630 32622 5682
rect 32622 5630 32674 5682
rect 32674 5630 32676 5682
rect 32620 5628 32676 5630
rect 32956 6578 33012 6580
rect 32956 6526 32958 6578
rect 32958 6526 33010 6578
rect 33010 6526 33012 6578
rect 32956 6524 33012 6526
rect 32844 5516 32900 5572
rect 32732 5180 32788 5236
rect 32620 5010 32676 5012
rect 32620 4958 32622 5010
rect 32622 4958 32674 5010
rect 32674 4958 32676 5010
rect 32620 4956 32676 4958
rect 32284 4284 32340 4340
rect 33516 7756 33572 7812
rect 33628 7420 33684 7476
rect 33964 6636 34020 6692
rect 32844 4508 32900 4564
rect 33180 5628 33236 5684
rect 33740 5234 33796 5236
rect 33740 5182 33742 5234
rect 33742 5182 33794 5234
rect 33794 5182 33796 5234
rect 33740 5180 33796 5182
rect 33404 4508 33460 4564
rect 32508 3330 32564 3332
rect 32508 3278 32510 3330
rect 32510 3278 32562 3330
rect 32562 3278 32564 3330
rect 32508 3276 32564 3278
rect 31164 2492 31220 2548
rect 32060 1484 32116 1540
rect 33628 4226 33684 4228
rect 33628 4174 33630 4226
rect 33630 4174 33682 4226
rect 33682 4174 33684 4226
rect 33628 4172 33684 4174
rect 34636 10108 34692 10164
rect 35420 13468 35476 13524
rect 35532 13692 35588 13748
rect 34972 13356 35028 13412
rect 34860 12124 34916 12180
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 13074 35252 13076
rect 35196 13022 35198 13074
rect 35198 13022 35250 13074
rect 35250 13022 35252 13074
rect 35196 13020 35252 13022
rect 35084 12290 35140 12292
rect 35084 12238 35086 12290
rect 35086 12238 35138 12290
rect 35138 12238 35140 12290
rect 35084 12236 35140 12238
rect 35308 12178 35364 12180
rect 35308 12126 35310 12178
rect 35310 12126 35362 12178
rect 35362 12126 35364 12178
rect 35308 12124 35364 12126
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34860 10892 34916 10948
rect 35532 10892 35588 10948
rect 34972 10780 35028 10836
rect 35980 16380 36036 16436
rect 37100 23042 37156 23044
rect 37100 22990 37102 23042
rect 37102 22990 37154 23042
rect 37154 22990 37156 23042
rect 37100 22988 37156 22990
rect 37324 21980 37380 22036
rect 36652 20690 36708 20692
rect 36652 20638 36654 20690
rect 36654 20638 36706 20690
rect 36706 20638 36708 20690
rect 36652 20636 36708 20638
rect 36540 20412 36596 20468
rect 36988 20188 37044 20244
rect 36764 19292 36820 19348
rect 36428 19180 36484 19236
rect 36652 18284 36708 18340
rect 36204 17052 36260 17108
rect 36540 17052 36596 17108
rect 36652 18060 36708 18116
rect 36316 16940 36372 16996
rect 36652 16828 36708 16884
rect 36204 16380 36260 16436
rect 36316 16098 36372 16100
rect 36316 16046 36318 16098
rect 36318 16046 36370 16098
rect 36370 16046 36372 16098
rect 36316 16044 36372 16046
rect 36316 15820 36372 15876
rect 36764 16380 36820 16436
rect 36876 18284 36932 18340
rect 36540 16156 36596 16212
rect 36540 15986 36596 15988
rect 36540 15934 36542 15986
rect 36542 15934 36594 15986
rect 36594 15934 36596 15986
rect 36540 15932 36596 15934
rect 36652 15874 36708 15876
rect 36652 15822 36654 15874
rect 36654 15822 36706 15874
rect 36706 15822 36708 15874
rect 36652 15820 36708 15822
rect 36652 15596 36708 15652
rect 36764 15484 36820 15540
rect 36316 15426 36372 15428
rect 36316 15374 36318 15426
rect 36318 15374 36370 15426
rect 36370 15374 36372 15426
rect 36316 15372 36372 15374
rect 36428 15260 36484 15316
rect 36204 14476 36260 14532
rect 35980 13858 36036 13860
rect 35980 13806 35982 13858
rect 35982 13806 36034 13858
rect 36034 13806 36036 13858
rect 35980 13804 36036 13806
rect 35868 13468 35924 13524
rect 35756 13020 35812 13076
rect 36092 12850 36148 12852
rect 36092 12798 36094 12850
rect 36094 12798 36146 12850
rect 36146 12798 36148 12850
rect 36092 12796 36148 12798
rect 36204 12572 36260 12628
rect 36316 13244 36372 13300
rect 35868 12236 35924 12292
rect 35756 12012 35812 12068
rect 36540 13692 36596 13748
rect 36652 13468 36708 13524
rect 36764 12850 36820 12852
rect 36764 12798 36766 12850
rect 36766 12798 36818 12850
rect 36818 12798 36820 12850
rect 36764 12796 36820 12798
rect 36428 12460 36484 12516
rect 36652 12402 36708 12404
rect 36652 12350 36654 12402
rect 36654 12350 36706 12402
rect 36706 12350 36708 12402
rect 36652 12348 36708 12350
rect 36764 12290 36820 12292
rect 36764 12238 36766 12290
rect 36766 12238 36818 12290
rect 36818 12238 36820 12290
rect 36764 12236 36820 12238
rect 36092 11564 36148 11620
rect 36092 11004 36148 11060
rect 36316 10892 36372 10948
rect 35980 10834 36036 10836
rect 35980 10782 35982 10834
rect 35982 10782 36034 10834
rect 36034 10782 36036 10834
rect 35980 10780 36036 10782
rect 34972 10610 35028 10612
rect 34972 10558 34974 10610
rect 34974 10558 35026 10610
rect 35026 10558 35028 10610
rect 34972 10556 35028 10558
rect 35308 10556 35364 10612
rect 35308 10332 35364 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34748 9042 34804 9044
rect 34748 8990 34750 9042
rect 34750 8990 34802 9042
rect 34802 8990 34804 9042
rect 34748 8988 34804 8990
rect 34860 8930 34916 8932
rect 34860 8878 34862 8930
rect 34862 8878 34914 8930
rect 34914 8878 34916 8930
rect 34860 8876 34916 8878
rect 34972 8764 35028 8820
rect 34860 7474 34916 7476
rect 34860 7422 34862 7474
rect 34862 7422 34914 7474
rect 34914 7422 34916 7474
rect 34860 7420 34916 7422
rect 35308 9938 35364 9940
rect 35308 9886 35310 9938
rect 35310 9886 35362 9938
rect 35362 9886 35364 9938
rect 35308 9884 35364 9886
rect 35980 10556 36036 10612
rect 35980 10108 36036 10164
rect 36092 10332 36148 10388
rect 35868 9996 35924 10052
rect 36764 11506 36820 11508
rect 36764 11454 36766 11506
rect 36766 11454 36818 11506
rect 36818 11454 36820 11506
rect 36764 11452 36820 11454
rect 36764 11228 36820 11284
rect 36652 11116 36708 11172
rect 36428 10332 36484 10388
rect 36540 10668 36596 10724
rect 36540 10220 36596 10276
rect 36764 10332 36820 10388
rect 36204 9772 36260 9828
rect 35532 9324 35588 9380
rect 35532 8930 35588 8932
rect 35532 8878 35534 8930
rect 35534 8878 35586 8930
rect 35586 8878 35588 8930
rect 35532 8876 35588 8878
rect 35420 8764 35476 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35980 9436 36036 9492
rect 36652 9154 36708 9156
rect 36652 9102 36654 9154
rect 36654 9102 36706 9154
rect 36706 9102 36708 9154
rect 36652 9100 36708 9102
rect 35644 8204 35700 8260
rect 35756 7980 35812 8036
rect 35532 7868 35588 7924
rect 35420 7756 35476 7812
rect 36428 8370 36484 8372
rect 36428 8318 36430 8370
rect 36430 8318 36482 8370
rect 36482 8318 36484 8370
rect 36428 8316 36484 8318
rect 36316 8204 36372 8260
rect 37212 19964 37268 20020
rect 37100 19906 37156 19908
rect 37100 19854 37102 19906
rect 37102 19854 37154 19906
rect 37154 19854 37156 19906
rect 37100 19852 37156 19854
rect 37100 18338 37156 18340
rect 37100 18286 37102 18338
rect 37102 18286 37154 18338
rect 37154 18286 37156 18338
rect 37100 18284 37156 18286
rect 37436 21868 37492 21924
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 37884 22370 37940 22372
rect 37884 22318 37886 22370
rect 37886 22318 37938 22370
rect 37938 22318 37940 22370
rect 37884 22316 37940 22318
rect 37884 21980 37940 22036
rect 37436 20802 37492 20804
rect 37436 20750 37438 20802
rect 37438 20750 37490 20802
rect 37490 20750 37492 20802
rect 37436 20748 37492 20750
rect 37996 20860 38052 20916
rect 37548 19628 37604 19684
rect 37436 18844 37492 18900
rect 37548 19180 37604 19236
rect 37212 17948 37268 18004
rect 37884 19964 37940 20020
rect 37996 20188 38052 20244
rect 37996 19740 38052 19796
rect 37772 18396 37828 18452
rect 37660 18338 37716 18340
rect 37660 18286 37662 18338
rect 37662 18286 37714 18338
rect 37714 18286 37716 18338
rect 37660 18284 37716 18286
rect 38108 19180 38164 19236
rect 38332 22428 38388 22484
rect 39452 23826 39508 23828
rect 39452 23774 39454 23826
rect 39454 23774 39506 23826
rect 39506 23774 39508 23826
rect 39452 23772 39508 23774
rect 38668 22428 38724 22484
rect 39004 22652 39060 22708
rect 38780 22316 38836 22372
rect 38892 22092 38948 22148
rect 38332 21644 38388 21700
rect 38444 21308 38500 21364
rect 38780 20972 38836 21028
rect 38444 19906 38500 19908
rect 38444 19854 38446 19906
rect 38446 19854 38498 19906
rect 38498 19854 38500 19906
rect 38444 19852 38500 19854
rect 38108 18956 38164 19012
rect 37100 17106 37156 17108
rect 37100 17054 37102 17106
rect 37102 17054 37154 17106
rect 37154 17054 37156 17106
rect 37100 17052 37156 17054
rect 37324 17106 37380 17108
rect 37324 17054 37326 17106
rect 37326 17054 37378 17106
rect 37378 17054 37380 17106
rect 37324 17052 37380 17054
rect 37324 16828 37380 16884
rect 37212 15932 37268 15988
rect 37212 15708 37268 15764
rect 37100 15426 37156 15428
rect 37100 15374 37102 15426
rect 37102 15374 37154 15426
rect 37154 15374 37156 15426
rect 37100 15372 37156 15374
rect 37100 14588 37156 14644
rect 36988 13522 37044 13524
rect 36988 13470 36990 13522
rect 36990 13470 37042 13522
rect 37042 13470 37044 13522
rect 36988 13468 37044 13470
rect 37436 16156 37492 16212
rect 37436 15596 37492 15652
rect 37436 15426 37492 15428
rect 37436 15374 37438 15426
rect 37438 15374 37490 15426
rect 37490 15374 37492 15426
rect 37436 15372 37492 15374
rect 37660 16044 37716 16100
rect 37772 15708 37828 15764
rect 38108 17612 38164 17668
rect 38108 17442 38164 17444
rect 38108 17390 38110 17442
rect 38110 17390 38162 17442
rect 38162 17390 38164 17442
rect 38108 17388 38164 17390
rect 38780 18844 38836 18900
rect 40236 23714 40292 23716
rect 40236 23662 40238 23714
rect 40238 23662 40290 23714
rect 40290 23662 40292 23714
rect 40236 23660 40292 23662
rect 40684 23548 40740 23604
rect 41244 23436 41300 23492
rect 39676 23266 39732 23268
rect 39676 23214 39678 23266
rect 39678 23214 39730 23266
rect 39730 23214 39732 23266
rect 39676 23212 39732 23214
rect 39228 23042 39284 23044
rect 39228 22990 39230 23042
rect 39230 22990 39282 23042
rect 39282 22990 39284 23042
rect 39228 22988 39284 22990
rect 39900 22540 39956 22596
rect 39676 21980 39732 22036
rect 39340 21756 39396 21812
rect 39340 21474 39396 21476
rect 39340 21422 39342 21474
rect 39342 21422 39394 21474
rect 39394 21422 39396 21474
rect 39340 21420 39396 21422
rect 39228 20578 39284 20580
rect 39228 20526 39230 20578
rect 39230 20526 39282 20578
rect 39282 20526 39284 20578
rect 39228 20524 39284 20526
rect 39340 20130 39396 20132
rect 39340 20078 39342 20130
rect 39342 20078 39394 20130
rect 39394 20078 39396 20130
rect 39340 20076 39396 20078
rect 39116 19852 39172 19908
rect 40012 21980 40068 22036
rect 39900 21868 39956 21924
rect 40572 22146 40628 22148
rect 40572 22094 40574 22146
rect 40574 22094 40626 22146
rect 40626 22094 40628 22146
rect 40572 22092 40628 22094
rect 40236 21644 40292 21700
rect 40460 21756 40516 21812
rect 39788 19516 39844 19572
rect 39676 19122 39732 19124
rect 39676 19070 39678 19122
rect 39678 19070 39730 19122
rect 39730 19070 39732 19122
rect 39676 19068 39732 19070
rect 39228 19010 39284 19012
rect 39228 18958 39230 19010
rect 39230 18958 39282 19010
rect 39282 18958 39284 19010
rect 39228 18956 39284 18958
rect 40012 20412 40068 20468
rect 39900 18844 39956 18900
rect 40012 18956 40068 19012
rect 39452 18450 39508 18452
rect 39452 18398 39454 18450
rect 39454 18398 39506 18450
rect 39506 18398 39508 18450
rect 39452 18396 39508 18398
rect 39900 18172 39956 18228
rect 38892 18060 38948 18116
rect 38444 17442 38500 17444
rect 38444 17390 38446 17442
rect 38446 17390 38498 17442
rect 38498 17390 38500 17442
rect 38444 17388 38500 17390
rect 38332 16994 38388 16996
rect 38332 16942 38334 16994
rect 38334 16942 38386 16994
rect 38386 16942 38388 16994
rect 38332 16940 38388 16942
rect 37996 16828 38052 16884
rect 37324 14588 37380 14644
rect 37212 13858 37268 13860
rect 37212 13806 37214 13858
rect 37214 13806 37266 13858
rect 37266 13806 37268 13858
rect 37212 13804 37268 13806
rect 38332 15426 38388 15428
rect 38332 15374 38334 15426
rect 38334 15374 38386 15426
rect 38386 15374 38388 15426
rect 38332 15372 38388 15374
rect 37436 14252 37492 14308
rect 37324 13244 37380 13300
rect 37548 13916 37604 13972
rect 37324 12796 37380 12852
rect 37100 11452 37156 11508
rect 37212 12460 37268 12516
rect 37100 10498 37156 10500
rect 37100 10446 37102 10498
rect 37102 10446 37154 10498
rect 37154 10446 37156 10498
rect 37100 10444 37156 10446
rect 37100 10220 37156 10276
rect 36876 8876 36932 8932
rect 36988 9436 37044 9492
rect 36316 8034 36372 8036
rect 36316 7982 36318 8034
rect 36318 7982 36370 8034
rect 36370 7982 36372 8034
rect 36316 7980 36372 7982
rect 36092 7868 36148 7924
rect 36764 7756 36820 7812
rect 35308 7362 35364 7364
rect 35308 7310 35310 7362
rect 35310 7310 35362 7362
rect 35362 7310 35364 7362
rect 35308 7308 35364 7310
rect 36316 7362 36372 7364
rect 36316 7310 36318 7362
rect 36318 7310 36370 7362
rect 36370 7310 36372 7362
rect 36316 7308 36372 7310
rect 35084 7250 35140 7252
rect 35084 7198 35086 7250
rect 35086 7198 35138 7250
rect 35138 7198 35140 7250
rect 35084 7196 35140 7198
rect 36540 7250 36596 7252
rect 36540 7198 36542 7250
rect 36542 7198 36594 7250
rect 36594 7198 36596 7250
rect 36540 7196 36596 7198
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 36764 7474 36820 7476
rect 36764 7422 36766 7474
rect 36766 7422 36818 7474
rect 36818 7422 36820 7474
rect 36764 7420 36820 7422
rect 35084 5964 35140 6020
rect 35980 6412 36036 6468
rect 36204 6300 36260 6356
rect 35980 5964 36036 6020
rect 35756 5794 35812 5796
rect 35756 5742 35758 5794
rect 35758 5742 35810 5794
rect 35810 5742 35812 5794
rect 35756 5740 35812 5742
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35756 5404 35812 5460
rect 35868 5346 35924 5348
rect 35868 5294 35870 5346
rect 35870 5294 35922 5346
rect 35922 5294 35924 5346
rect 35868 5292 35924 5294
rect 34524 5068 34580 5124
rect 34972 4508 35028 4564
rect 36204 5516 36260 5572
rect 36092 5122 36148 5124
rect 36092 5070 36094 5122
rect 36094 5070 36146 5122
rect 36146 5070 36148 5122
rect 36092 5068 36148 5070
rect 36316 5122 36372 5124
rect 36316 5070 36318 5122
rect 36318 5070 36370 5122
rect 36370 5070 36372 5122
rect 36316 5068 36372 5070
rect 36428 4338 36484 4340
rect 36428 4286 36430 4338
rect 36430 4286 36482 4338
rect 36482 4286 36484 4338
rect 36428 4284 36484 4286
rect 34300 4060 34356 4116
rect 35532 4060 35588 4116
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35756 3778 35812 3780
rect 35756 3726 35758 3778
rect 35758 3726 35810 3778
rect 35810 3726 35812 3778
rect 35756 3724 35812 3726
rect 35868 3666 35924 3668
rect 35868 3614 35870 3666
rect 35870 3614 35922 3666
rect 35922 3614 35924 3666
rect 35868 3612 35924 3614
rect 34524 1484 34580 1540
rect 34748 3388 34804 3444
rect 35420 3164 35476 3220
rect 36988 7756 37044 7812
rect 36876 5964 36932 6020
rect 38108 14306 38164 14308
rect 38108 14254 38110 14306
rect 38110 14254 38162 14306
rect 38162 14254 38164 14306
rect 38108 14252 38164 14254
rect 38668 17106 38724 17108
rect 38668 17054 38670 17106
rect 38670 17054 38722 17106
rect 38722 17054 38724 17106
rect 38668 17052 38724 17054
rect 38556 15372 38612 15428
rect 38668 16380 38724 16436
rect 39004 17388 39060 17444
rect 39116 16098 39172 16100
rect 39116 16046 39118 16098
rect 39118 16046 39170 16098
rect 39170 16046 39172 16098
rect 39116 16044 39172 16046
rect 38892 15932 38948 15988
rect 38780 15314 38836 15316
rect 38780 15262 38782 15314
rect 38782 15262 38834 15314
rect 38834 15262 38836 15314
rect 38780 15260 38836 15262
rect 39340 17442 39396 17444
rect 39340 17390 39342 17442
rect 39342 17390 39394 17442
rect 39394 17390 39396 17442
rect 39340 17388 39396 17390
rect 40348 19906 40404 19908
rect 40348 19854 40350 19906
rect 40350 19854 40402 19906
rect 40402 19854 40404 19906
rect 40348 19852 40404 19854
rect 40460 19740 40516 19796
rect 41020 21868 41076 21924
rect 43148 24444 43204 24500
rect 42476 24108 42532 24164
rect 41580 23100 41636 23156
rect 41468 23042 41524 23044
rect 41468 22990 41470 23042
rect 41470 22990 41522 23042
rect 41522 22990 41524 23042
rect 41468 22988 41524 22990
rect 41356 22540 41412 22596
rect 41692 21868 41748 21924
rect 42028 23266 42084 23268
rect 42028 23214 42030 23266
rect 42030 23214 42082 23266
rect 42082 23214 42084 23266
rect 42028 23212 42084 23214
rect 42364 23212 42420 23268
rect 42140 22428 42196 22484
rect 41804 21756 41860 21812
rect 40684 19292 40740 19348
rect 41916 21420 41972 21476
rect 41580 20860 41636 20916
rect 41468 19906 41524 19908
rect 41468 19854 41470 19906
rect 41470 19854 41522 19906
rect 41522 19854 41524 19906
rect 41468 19852 41524 19854
rect 41356 19404 41412 19460
rect 41356 19180 41412 19236
rect 40012 17164 40068 17220
rect 40124 17724 40180 17780
rect 39340 16882 39396 16884
rect 39340 16830 39342 16882
rect 39342 16830 39394 16882
rect 39394 16830 39396 16882
rect 39340 16828 39396 16830
rect 39788 16940 39844 16996
rect 39676 16882 39732 16884
rect 39676 16830 39678 16882
rect 39678 16830 39730 16882
rect 39730 16830 39732 16882
rect 39676 16828 39732 16830
rect 39564 16210 39620 16212
rect 39564 16158 39566 16210
rect 39566 16158 39618 16210
rect 39618 16158 39620 16210
rect 39564 16156 39620 16158
rect 39340 16044 39396 16100
rect 39452 15932 39508 15988
rect 39900 16380 39956 16436
rect 39900 15820 39956 15876
rect 39564 15426 39620 15428
rect 39564 15374 39566 15426
rect 39566 15374 39618 15426
rect 39618 15374 39620 15426
rect 39564 15372 39620 15374
rect 38892 14812 38948 14868
rect 38444 14140 38500 14196
rect 37772 14028 37828 14084
rect 37660 13020 37716 13076
rect 37772 13804 37828 13860
rect 38332 13858 38388 13860
rect 38332 13806 38334 13858
rect 38334 13806 38386 13858
rect 38386 13806 38388 13858
rect 38332 13804 38388 13806
rect 38220 13692 38276 13748
rect 38108 13522 38164 13524
rect 38108 13470 38110 13522
rect 38110 13470 38162 13522
rect 38162 13470 38164 13522
rect 38108 13468 38164 13470
rect 39116 14418 39172 14420
rect 39116 14366 39118 14418
rect 39118 14366 39170 14418
rect 39170 14366 39172 14418
rect 39116 14364 39172 14366
rect 39900 14588 39956 14644
rect 40012 15708 40068 15764
rect 39564 14418 39620 14420
rect 39564 14366 39566 14418
rect 39566 14366 39618 14418
rect 39618 14366 39620 14418
rect 39564 14364 39620 14366
rect 39900 14418 39956 14420
rect 39900 14366 39902 14418
rect 39902 14366 39954 14418
rect 39954 14366 39956 14418
rect 39900 14364 39956 14366
rect 39564 13970 39620 13972
rect 39564 13918 39566 13970
rect 39566 13918 39618 13970
rect 39618 13918 39620 13970
rect 39564 13916 39620 13918
rect 39676 13804 39732 13860
rect 39340 13356 39396 13412
rect 39116 13020 39172 13076
rect 38556 12908 38612 12964
rect 37660 12850 37716 12852
rect 37660 12798 37662 12850
rect 37662 12798 37714 12850
rect 37714 12798 37716 12850
rect 37660 12796 37716 12798
rect 38108 12796 38164 12852
rect 37772 12684 37828 12740
rect 37436 11788 37492 11844
rect 37548 11676 37604 11732
rect 37660 12124 37716 12180
rect 37324 11452 37380 11508
rect 37772 11452 37828 11508
rect 37436 11170 37492 11172
rect 37436 11118 37438 11170
rect 37438 11118 37490 11170
rect 37490 11118 37492 11170
rect 37436 11116 37492 11118
rect 37660 11282 37716 11284
rect 37660 11230 37662 11282
rect 37662 11230 37714 11282
rect 37714 11230 37716 11282
rect 37660 11228 37716 11230
rect 38668 12962 38724 12964
rect 38668 12910 38670 12962
rect 38670 12910 38722 12962
rect 38722 12910 38724 12962
rect 38668 12908 38724 12910
rect 38780 12738 38836 12740
rect 38780 12686 38782 12738
rect 38782 12686 38834 12738
rect 38834 12686 38836 12738
rect 38780 12684 38836 12686
rect 38444 12402 38500 12404
rect 38444 12350 38446 12402
rect 38446 12350 38498 12402
rect 38498 12350 38500 12402
rect 38444 12348 38500 12350
rect 38668 12290 38724 12292
rect 38668 12238 38670 12290
rect 38670 12238 38722 12290
rect 38722 12238 38724 12290
rect 38668 12236 38724 12238
rect 38108 11954 38164 11956
rect 38108 11902 38110 11954
rect 38110 11902 38162 11954
rect 38162 11902 38164 11954
rect 38108 11900 38164 11902
rect 38556 12012 38612 12068
rect 37884 11228 37940 11284
rect 38444 11282 38500 11284
rect 38444 11230 38446 11282
rect 38446 11230 38498 11282
rect 38498 11230 38500 11282
rect 38444 11228 38500 11230
rect 38780 12012 38836 12068
rect 39004 12850 39060 12852
rect 39004 12798 39006 12850
rect 39006 12798 39058 12850
rect 39058 12798 39060 12850
rect 39004 12796 39060 12798
rect 38444 11004 38500 11060
rect 38668 11452 38724 11508
rect 37436 10610 37492 10612
rect 37436 10558 37438 10610
rect 37438 10558 37490 10610
rect 37490 10558 37492 10610
rect 37436 10556 37492 10558
rect 37660 10610 37716 10612
rect 37660 10558 37662 10610
rect 37662 10558 37714 10610
rect 37714 10558 37716 10610
rect 37660 10556 37716 10558
rect 38444 10780 38500 10836
rect 38892 11004 38948 11060
rect 38220 10444 38276 10500
rect 37772 9996 37828 10052
rect 37548 9826 37604 9828
rect 37548 9774 37550 9826
rect 37550 9774 37602 9826
rect 37602 9774 37604 9826
rect 37548 9772 37604 9774
rect 37884 9884 37940 9940
rect 37324 9436 37380 9492
rect 37324 8818 37380 8820
rect 37324 8766 37326 8818
rect 37326 8766 37378 8818
rect 37378 8766 37380 8818
rect 37324 8764 37380 8766
rect 37660 9436 37716 9492
rect 37996 9042 38052 9044
rect 37996 8990 37998 9042
rect 37998 8990 38050 9042
rect 38050 8990 38052 9042
rect 37996 8988 38052 8990
rect 37660 8652 37716 8708
rect 38108 8652 38164 8708
rect 38556 9826 38612 9828
rect 38556 9774 38558 9826
rect 38558 9774 38610 9826
rect 38610 9774 38612 9826
rect 38556 9772 38612 9774
rect 38780 9772 38836 9828
rect 38444 8652 38500 8708
rect 37772 8146 37828 8148
rect 37772 8094 37774 8146
rect 37774 8094 37826 8146
rect 37826 8094 37828 8146
rect 37772 8092 37828 8094
rect 37324 7756 37380 7812
rect 37884 7980 37940 8036
rect 38668 8428 38724 8484
rect 38108 8204 38164 8260
rect 37212 7084 37268 7140
rect 38332 8204 38388 8260
rect 37212 6076 37268 6132
rect 38332 7756 38388 7812
rect 38220 6130 38276 6132
rect 38220 6078 38222 6130
rect 38222 6078 38274 6130
rect 38274 6078 38276 6130
rect 38220 6076 38276 6078
rect 37772 6018 37828 6020
rect 37772 5966 37774 6018
rect 37774 5966 37826 6018
rect 37826 5966 37828 6018
rect 37772 5964 37828 5966
rect 36988 5068 37044 5124
rect 37100 5180 37156 5236
rect 37436 5794 37492 5796
rect 37436 5742 37438 5794
rect 37438 5742 37490 5794
rect 37490 5742 37492 5794
rect 37436 5740 37492 5742
rect 37772 5740 37828 5796
rect 37660 5292 37716 5348
rect 37212 3276 37268 3332
rect 37436 4732 37492 4788
rect 36540 3052 36596 3108
rect 35420 2828 35476 2884
rect 35308 2604 35364 2660
rect 34748 2380 34804 2436
rect 36092 2044 36148 2100
rect 37772 3724 37828 3780
rect 38444 6690 38500 6692
rect 38444 6638 38446 6690
rect 38446 6638 38498 6690
rect 38498 6638 38500 6690
rect 38444 6636 38500 6638
rect 38556 5292 38612 5348
rect 39676 12962 39732 12964
rect 39676 12910 39678 12962
rect 39678 12910 39730 12962
rect 39730 12910 39732 12962
rect 39676 12908 39732 12910
rect 40012 13356 40068 13412
rect 39900 12850 39956 12852
rect 39900 12798 39902 12850
rect 39902 12798 39954 12850
rect 39954 12798 39956 12850
rect 39900 12796 39956 12798
rect 39452 12348 39508 12404
rect 39116 11228 39172 11284
rect 39452 11340 39508 11396
rect 39564 10780 39620 10836
rect 39004 9436 39060 9492
rect 39228 9436 39284 9492
rect 39228 9212 39284 9268
rect 39564 9884 39620 9940
rect 39788 12684 39844 12740
rect 40012 11564 40068 11620
rect 39788 11394 39844 11396
rect 39788 11342 39790 11394
rect 39790 11342 39842 11394
rect 39842 11342 39844 11394
rect 39788 11340 39844 11342
rect 39788 10108 39844 10164
rect 40684 19010 40740 19012
rect 40684 18958 40686 19010
rect 40686 18958 40738 19010
rect 40738 18958 40740 19010
rect 40684 18956 40740 18958
rect 40460 18508 40516 18564
rect 40684 18396 40740 18452
rect 40460 17836 40516 17892
rect 40460 17276 40516 17332
rect 40572 17164 40628 17220
rect 40796 18338 40852 18340
rect 40796 18286 40798 18338
rect 40798 18286 40850 18338
rect 40850 18286 40852 18338
rect 40796 18284 40852 18286
rect 40572 16994 40628 16996
rect 40572 16942 40574 16994
rect 40574 16942 40626 16994
rect 40626 16942 40628 16994
rect 40572 16940 40628 16942
rect 40460 16882 40516 16884
rect 40460 16830 40462 16882
rect 40462 16830 40514 16882
rect 40514 16830 40516 16882
rect 40460 16828 40516 16830
rect 40348 16492 40404 16548
rect 40572 15986 40628 15988
rect 40572 15934 40574 15986
rect 40574 15934 40626 15986
rect 40626 15934 40628 15986
rect 40572 15932 40628 15934
rect 40348 15708 40404 15764
rect 40460 15596 40516 15652
rect 40572 15708 40628 15764
rect 40236 15484 40292 15540
rect 40236 15314 40292 15316
rect 40236 15262 40238 15314
rect 40238 15262 40290 15314
rect 40290 15262 40292 15314
rect 40236 15260 40292 15262
rect 40236 14588 40292 14644
rect 41020 16604 41076 16660
rect 41020 15874 41076 15876
rect 41020 15822 41022 15874
rect 41022 15822 41074 15874
rect 41074 15822 41076 15874
rect 41020 15820 41076 15822
rect 40684 15260 40740 15316
rect 40684 14418 40740 14420
rect 40684 14366 40686 14418
rect 40686 14366 40738 14418
rect 40738 14366 40740 14418
rect 40684 14364 40740 14366
rect 40572 13916 40628 13972
rect 40684 14140 40740 14196
rect 40572 13746 40628 13748
rect 40572 13694 40574 13746
rect 40574 13694 40626 13746
rect 40626 13694 40628 13746
rect 40572 13692 40628 13694
rect 40684 13580 40740 13636
rect 40572 12962 40628 12964
rect 40572 12910 40574 12962
rect 40574 12910 40626 12962
rect 40626 12910 40628 12962
rect 40572 12908 40628 12910
rect 40684 12738 40740 12740
rect 40684 12686 40686 12738
rect 40686 12686 40738 12738
rect 40738 12686 40740 12738
rect 40684 12684 40740 12686
rect 40572 12572 40628 12628
rect 40460 12124 40516 12180
rect 40236 11452 40292 11508
rect 40236 11004 40292 11060
rect 40460 11618 40516 11620
rect 40460 11566 40462 11618
rect 40462 11566 40514 11618
rect 40514 11566 40516 11618
rect 40460 11564 40516 11566
rect 40460 11282 40516 11284
rect 40460 11230 40462 11282
rect 40462 11230 40514 11282
rect 40514 11230 40516 11282
rect 40460 11228 40516 11230
rect 40572 11116 40628 11172
rect 41020 12348 41076 12404
rect 40908 12236 40964 12292
rect 40348 10892 40404 10948
rect 41244 17948 41300 18004
rect 41468 18284 41524 18340
rect 41356 17388 41412 17444
rect 41244 17052 41300 17108
rect 42028 20914 42084 20916
rect 42028 20862 42030 20914
rect 42030 20862 42082 20914
rect 42082 20862 42084 20914
rect 42028 20860 42084 20862
rect 41804 18172 41860 18228
rect 42028 19346 42084 19348
rect 42028 19294 42030 19346
rect 42030 19294 42082 19346
rect 42082 19294 42084 19346
rect 42028 19292 42084 19294
rect 42028 18338 42084 18340
rect 42028 18286 42030 18338
rect 42030 18286 42082 18338
rect 42082 18286 42084 18338
rect 42028 18284 42084 18286
rect 41916 18060 41972 18116
rect 41692 17836 41748 17892
rect 41916 17836 41972 17892
rect 41580 17724 41636 17780
rect 41916 17276 41972 17332
rect 41468 16044 41524 16100
rect 41580 17164 41636 17220
rect 41692 16604 41748 16660
rect 41804 16716 41860 16772
rect 41916 16380 41972 16436
rect 41804 16098 41860 16100
rect 41804 16046 41806 16098
rect 41806 16046 41858 16098
rect 41858 16046 41860 16098
rect 41804 16044 41860 16046
rect 41468 15874 41524 15876
rect 41468 15822 41470 15874
rect 41470 15822 41522 15874
rect 41522 15822 41524 15874
rect 41468 15820 41524 15822
rect 41692 15260 41748 15316
rect 41468 15148 41524 15204
rect 41804 15148 41860 15204
rect 41356 14252 41412 14308
rect 41916 14476 41972 14532
rect 41580 14140 41636 14196
rect 41692 14306 41748 14308
rect 41692 14254 41694 14306
rect 41694 14254 41746 14306
rect 41746 14254 41748 14306
rect 41692 14252 41748 14254
rect 41692 13970 41748 13972
rect 41692 13918 41694 13970
rect 41694 13918 41746 13970
rect 41746 13918 41748 13970
rect 41692 13916 41748 13918
rect 41244 13692 41300 13748
rect 41468 12962 41524 12964
rect 41468 12910 41470 12962
rect 41470 12910 41522 12962
rect 41522 12910 41524 12962
rect 41468 12908 41524 12910
rect 41244 11282 41300 11284
rect 41244 11230 41246 11282
rect 41246 11230 41298 11282
rect 41298 11230 41300 11282
rect 41244 11228 41300 11230
rect 40460 10444 40516 10500
rect 40348 9996 40404 10052
rect 39788 9548 39844 9604
rect 39452 9266 39508 9268
rect 39452 9214 39454 9266
rect 39454 9214 39506 9266
rect 39506 9214 39508 9266
rect 39452 9212 39508 9214
rect 39340 8764 39396 8820
rect 39004 8428 39060 8484
rect 39340 8540 39396 8596
rect 39004 7980 39060 8036
rect 38892 7756 38948 7812
rect 39116 7698 39172 7700
rect 39116 7646 39118 7698
rect 39118 7646 39170 7698
rect 39170 7646 39172 7698
rect 39116 7644 39172 7646
rect 39676 9436 39732 9492
rect 39900 9436 39956 9492
rect 39788 9324 39844 9380
rect 39676 8988 39732 9044
rect 39564 8316 39620 8372
rect 39676 8092 39732 8148
rect 39788 8034 39844 8036
rect 39788 7982 39790 8034
rect 39790 7982 39842 8034
rect 39842 7982 39844 8034
rect 39788 7980 39844 7982
rect 39228 6860 39284 6916
rect 38780 6412 38836 6468
rect 38892 5794 38948 5796
rect 38892 5742 38894 5794
rect 38894 5742 38946 5794
rect 38946 5742 38948 5794
rect 38892 5740 38948 5742
rect 38332 4620 38388 4676
rect 38892 4732 38948 4788
rect 38332 3500 38388 3556
rect 38108 3442 38164 3444
rect 38108 3390 38110 3442
rect 38110 3390 38162 3442
rect 38162 3390 38164 3442
rect 38108 3388 38164 3390
rect 38444 2828 38500 2884
rect 38444 2044 38500 2100
rect 38668 1596 38724 1652
rect 38780 4396 38836 4452
rect 39116 5404 39172 5460
rect 39900 7644 39956 7700
rect 40348 9772 40404 9828
rect 40572 9714 40628 9716
rect 40572 9662 40574 9714
rect 40574 9662 40626 9714
rect 40626 9662 40628 9714
rect 40572 9660 40628 9662
rect 40572 9154 40628 9156
rect 40572 9102 40574 9154
rect 40574 9102 40626 9154
rect 40626 9102 40628 9154
rect 40572 9100 40628 9102
rect 40460 8988 40516 9044
rect 40796 9996 40852 10052
rect 40908 10108 40964 10164
rect 40796 9772 40852 9828
rect 40796 8988 40852 9044
rect 40908 9548 40964 9604
rect 40348 8652 40404 8708
rect 40236 7980 40292 8036
rect 40348 8316 40404 8372
rect 40124 7756 40180 7812
rect 40684 8370 40740 8372
rect 40684 8318 40686 8370
rect 40686 8318 40738 8370
rect 40738 8318 40740 8370
rect 40684 8316 40740 8318
rect 40684 7420 40740 7476
rect 40684 7084 40740 7140
rect 40572 6860 40628 6916
rect 40796 6748 40852 6804
rect 39900 6578 39956 6580
rect 39900 6526 39902 6578
rect 39902 6526 39954 6578
rect 39954 6526 39956 6578
rect 39900 6524 39956 6526
rect 41468 9996 41524 10052
rect 41356 9602 41412 9604
rect 41356 9550 41358 9602
rect 41358 9550 41410 9602
rect 41410 9550 41412 9602
rect 41356 9548 41412 9550
rect 41692 13244 41748 13300
rect 41692 12572 41748 12628
rect 41916 13356 41972 13412
rect 41692 12402 41748 12404
rect 41692 12350 41694 12402
rect 41694 12350 41746 12402
rect 41746 12350 41748 12402
rect 41692 12348 41748 12350
rect 42252 21868 42308 21924
rect 42364 20860 42420 20916
rect 42812 23884 42868 23940
rect 42476 17948 42532 18004
rect 42588 22316 42644 22372
rect 42252 17612 42308 17668
rect 42140 13244 42196 13300
rect 42364 14028 42420 14084
rect 42252 13020 42308 13076
rect 42028 12684 42084 12740
rect 41916 12012 41972 12068
rect 41692 10834 41748 10836
rect 41692 10782 41694 10834
rect 41694 10782 41746 10834
rect 41746 10782 41748 10834
rect 41692 10780 41748 10782
rect 42140 11228 42196 11284
rect 41692 10386 41748 10388
rect 41692 10334 41694 10386
rect 41694 10334 41746 10386
rect 41746 10334 41748 10386
rect 41692 10332 41748 10334
rect 41692 9714 41748 9716
rect 41692 9662 41694 9714
rect 41694 9662 41746 9714
rect 41746 9662 41748 9714
rect 41692 9660 41748 9662
rect 41916 9772 41972 9828
rect 41020 8540 41076 8596
rect 41020 8146 41076 8148
rect 41020 8094 41022 8146
rect 41022 8094 41074 8146
rect 41074 8094 41076 8146
rect 41020 8092 41076 8094
rect 41356 8764 41412 8820
rect 41244 8652 41300 8708
rect 41244 7644 41300 7700
rect 41804 9212 41860 9268
rect 41692 9154 41748 9156
rect 41692 9102 41694 9154
rect 41694 9102 41746 9154
rect 41746 9102 41748 9154
rect 41692 9100 41748 9102
rect 41356 7196 41412 7252
rect 41468 8092 41524 8148
rect 41244 6466 41300 6468
rect 41244 6414 41246 6466
rect 41246 6414 41298 6466
rect 41298 6414 41300 6466
rect 41244 6412 41300 6414
rect 40124 6018 40180 6020
rect 40124 5966 40126 6018
rect 40126 5966 40178 6018
rect 40178 5966 40180 6018
rect 40124 5964 40180 5966
rect 41132 5964 41188 6020
rect 39788 4956 39844 5012
rect 40236 4844 40292 4900
rect 40124 4450 40180 4452
rect 40124 4398 40126 4450
rect 40126 4398 40178 4450
rect 40178 4398 40180 4450
rect 40124 4396 40180 4398
rect 39676 4172 39732 4228
rect 39004 3724 39060 3780
rect 39788 3724 39844 3780
rect 39116 3554 39172 3556
rect 39116 3502 39118 3554
rect 39118 3502 39170 3554
rect 39170 3502 39172 3554
rect 39116 3500 39172 3502
rect 39564 3554 39620 3556
rect 39564 3502 39566 3554
rect 39566 3502 39618 3554
rect 39618 3502 39620 3554
rect 39564 3500 39620 3502
rect 39340 3442 39396 3444
rect 39340 3390 39342 3442
rect 39342 3390 39394 3442
rect 39394 3390 39396 3442
rect 39340 3388 39396 3390
rect 40124 3330 40180 3332
rect 40124 3278 40126 3330
rect 40126 3278 40178 3330
rect 40178 3278 40180 3330
rect 40124 3276 40180 3278
rect 40684 4844 40740 4900
rect 40908 3554 40964 3556
rect 40908 3502 40910 3554
rect 40910 3502 40962 3554
rect 40962 3502 40964 3554
rect 40908 3500 40964 3502
rect 41692 8146 41748 8148
rect 41692 8094 41694 8146
rect 41694 8094 41746 8146
rect 41746 8094 41748 8146
rect 41692 8092 41748 8094
rect 41580 7980 41636 8036
rect 41804 7868 41860 7924
rect 42140 8876 42196 8932
rect 41916 7756 41972 7812
rect 41692 7698 41748 7700
rect 41692 7646 41694 7698
rect 41694 7646 41746 7698
rect 41746 7646 41748 7698
rect 41692 7644 41748 7646
rect 41916 7308 41972 7364
rect 41692 7250 41748 7252
rect 41692 7198 41694 7250
rect 41694 7198 41746 7250
rect 41746 7198 41748 7250
rect 41692 7196 41748 7198
rect 41804 6860 41860 6916
rect 42028 7084 42084 7140
rect 41804 6188 41860 6244
rect 41692 6130 41748 6132
rect 41692 6078 41694 6130
rect 41694 6078 41746 6130
rect 41746 6078 41748 6130
rect 41692 6076 41748 6078
rect 41804 5346 41860 5348
rect 41804 5294 41806 5346
rect 41806 5294 41858 5346
rect 41858 5294 41860 5346
rect 41804 5292 41860 5294
rect 41244 5068 41300 5124
rect 41580 5180 41636 5236
rect 41916 5122 41972 5124
rect 41916 5070 41918 5122
rect 41918 5070 41970 5122
rect 41970 5070 41972 5122
rect 41916 5068 41972 5070
rect 41804 5010 41860 5012
rect 41804 4958 41806 5010
rect 41806 4958 41858 5010
rect 41858 4958 41860 5010
rect 41804 4956 41860 4958
rect 41804 4338 41860 4340
rect 41804 4286 41806 4338
rect 41806 4286 41858 4338
rect 41858 4286 41860 4338
rect 41804 4284 41860 4286
rect 41580 3724 41636 3780
rect 41356 3554 41412 3556
rect 41356 3502 41358 3554
rect 41358 3502 41410 3554
rect 41410 3502 41412 3554
rect 41356 3500 41412 3502
rect 42140 6076 42196 6132
rect 42252 4508 42308 4564
rect 42700 22092 42756 22148
rect 42476 8428 42532 8484
rect 42588 13692 42644 13748
rect 42364 3724 42420 3780
rect 38780 2940 38836 2996
rect 41468 3276 41524 3332
rect 42588 2492 42644 2548
rect 42812 13020 42868 13076
rect 42924 23772 42980 23828
rect 42700 1484 42756 1540
rect 42812 6524 42868 6580
rect 42924 4732 42980 4788
rect 43036 22988 43092 23044
rect 43148 16940 43204 16996
rect 43260 10220 43316 10276
rect 43372 16828 43428 16884
rect 43036 2828 43092 2884
rect 43372 2604 43428 2660
<< metal3 >>
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 18386 39004 18396 39060
rect 18452 39004 21980 39060
rect 22036 39004 22046 39060
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 30034 27020 30044 27076
rect 30100 27020 36316 27076
rect 36372 27020 36382 27076
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 33058 25228 33068 25284
rect 33124 25228 43260 25284
rect 43316 25228 43326 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14354 24780 14364 24836
rect 14420 24780 38444 24836
rect 38500 24780 38510 24836
rect 30482 24668 30492 24724
rect 30548 24668 35756 24724
rect 35812 24668 35822 24724
rect 27010 24556 27020 24612
rect 27076 24556 30604 24612
rect 30660 24556 35980 24612
rect 36036 24556 36046 24612
rect 31892 24444 43148 24500
rect 43204 24444 43214 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 18386 23996 18396 24052
rect 18452 23996 28028 24052
rect 28084 23996 28094 24052
rect 31892 23940 31948 24444
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 25218 23884 25228 23940
rect 25284 23884 31948 23940
rect 33964 24108 42476 24164
rect 42532 24108 42542 24164
rect 33964 23828 34020 24108
rect 35746 23996 35756 24052
rect 35812 23996 36876 24052
rect 36932 23996 37548 24052
rect 37604 23996 37614 24052
rect 34178 23884 34188 23940
rect 34244 23884 42812 23940
rect 42868 23884 42878 23940
rect 24770 23772 24780 23828
rect 24836 23772 34020 23828
rect 39442 23772 39452 23828
rect 39508 23772 42924 23828
rect 42980 23772 42990 23828
rect 32610 23660 32620 23716
rect 32676 23660 33292 23716
rect 33348 23660 33358 23716
rect 35298 23660 35308 23716
rect 35364 23660 39340 23716
rect 39396 23660 39406 23716
rect 40114 23660 40124 23716
rect 40180 23660 40236 23716
rect 40292 23660 40302 23716
rect 26002 23548 26012 23604
rect 26068 23548 30492 23604
rect 30548 23548 30558 23604
rect 32498 23548 32508 23604
rect 32564 23548 36932 23604
rect 39890 23548 39900 23604
rect 39956 23548 40684 23604
rect 40740 23548 40750 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 36876 23492 36932 23548
rect 36876 23436 41244 23492
rect 41300 23436 41310 23492
rect 28690 23212 28700 23268
rect 28756 23212 31724 23268
rect 31780 23212 31790 23268
rect 32162 23212 32172 23268
rect 32228 23212 32508 23268
rect 32564 23212 33404 23268
rect 33460 23212 39676 23268
rect 39732 23212 39742 23268
rect 39900 23212 42028 23268
rect 42084 23212 42364 23268
rect 42420 23212 42430 23268
rect 39900 23156 39956 23212
rect 26450 23100 26460 23156
rect 26516 23100 29708 23156
rect 29764 23100 30828 23156
rect 30884 23100 30894 23156
rect 31826 23100 31836 23156
rect 31892 23100 35084 23156
rect 35140 23100 35150 23156
rect 37650 23100 37660 23156
rect 37716 23100 39956 23156
rect 40012 23100 41580 23156
rect 41636 23100 41646 23156
rect 40012 23044 40068 23100
rect 25554 22988 25564 23044
rect 25620 22988 26572 23044
rect 26628 22988 32620 23044
rect 32676 22988 33516 23044
rect 33572 22988 33852 23044
rect 33908 22988 34188 23044
rect 34244 22988 37100 23044
rect 37156 22988 37166 23044
rect 39218 22988 39228 23044
rect 39284 22988 40012 23044
rect 40068 22988 40078 23044
rect 41458 22988 41468 23044
rect 41524 22988 43036 23044
rect 43092 22988 43102 23044
rect 28578 22876 28588 22932
rect 28644 22876 28812 22932
rect 28868 22876 30044 22932
rect 30100 22876 30110 22932
rect 30594 22876 30604 22932
rect 30660 22876 33964 22932
rect 34020 22876 34030 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 29922 22652 29932 22708
rect 29988 22652 31388 22708
rect 31444 22652 31948 22708
rect 36418 22652 36428 22708
rect 36484 22652 39004 22708
rect 39060 22652 39070 22708
rect 31892 22596 31948 22652
rect 28242 22540 28252 22596
rect 28308 22540 30492 22596
rect 30548 22540 30558 22596
rect 30706 22540 30716 22596
rect 30772 22540 31500 22596
rect 31556 22540 31566 22596
rect 31892 22540 36540 22596
rect 36596 22540 36606 22596
rect 39890 22540 39900 22596
rect 39956 22540 41356 22596
rect 41412 22540 41422 22596
rect 23314 22428 23324 22484
rect 23380 22428 25564 22484
rect 25620 22428 25630 22484
rect 28802 22428 28812 22484
rect 28868 22428 29484 22484
rect 29540 22428 38332 22484
rect 38388 22428 38398 22484
rect 38658 22428 38668 22484
rect 38724 22428 42140 22484
rect 42196 22428 42206 22484
rect 3378 22316 3388 22372
rect 3444 22316 8428 22372
rect 8484 22316 8494 22372
rect 29474 22316 29484 22372
rect 29540 22316 30044 22372
rect 30100 22316 30110 22372
rect 30482 22316 30492 22372
rect 30548 22316 32508 22372
rect 32564 22316 32574 22372
rect 35074 22316 35084 22372
rect 35140 22316 37884 22372
rect 37940 22316 37950 22372
rect 38770 22316 38780 22372
rect 38836 22316 42588 22372
rect 42644 22316 42654 22372
rect 25554 22204 25564 22260
rect 25620 22204 27804 22260
rect 27860 22204 30268 22260
rect 30324 22204 30604 22260
rect 30660 22204 30670 22260
rect 31826 22204 31836 22260
rect 31892 22204 40684 22260
rect 40740 22204 40750 22260
rect 18610 22092 18620 22148
rect 18676 22092 24780 22148
rect 24836 22092 24846 22148
rect 26898 22092 26908 22148
rect 26964 22092 30604 22148
rect 30660 22092 30670 22148
rect 31266 22092 31276 22148
rect 31332 22092 33740 22148
rect 33796 22092 34972 22148
rect 35028 22092 35532 22148
rect 35588 22092 38892 22148
rect 38948 22092 38958 22148
rect 40562 22092 40572 22148
rect 40628 22092 42700 22148
rect 42756 22092 42766 22148
rect 0 22036 800 22064
rect 43200 22036 44000 22064
rect 0 21980 1820 22036
rect 1876 21980 1886 22036
rect 26226 21980 26236 22036
rect 26292 21980 34300 22036
rect 34356 21980 34366 22036
rect 34514 21980 34524 22036
rect 34580 21980 35084 22036
rect 35140 21980 35868 22036
rect 35924 21980 37324 22036
rect 37380 21980 37390 22036
rect 37874 21980 37884 22036
rect 37940 21980 39676 22036
rect 39732 21980 39742 22036
rect 40002 21980 40012 22036
rect 40068 21980 44000 22036
rect 0 21952 800 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 43200 21952 44000 21980
rect 21634 21868 21644 21924
rect 21700 21868 26908 21924
rect 26964 21868 26974 21924
rect 29334 21868 29372 21924
rect 29428 21868 29438 21924
rect 30930 21868 30940 21924
rect 30996 21868 35756 21924
rect 35812 21868 35822 21924
rect 37426 21868 37436 21924
rect 37492 21868 39900 21924
rect 39956 21868 39966 21924
rect 40674 21868 40684 21924
rect 40740 21868 41020 21924
rect 41076 21868 41086 21924
rect 41682 21868 41692 21924
rect 41748 21868 42252 21924
rect 42308 21868 42318 21924
rect 28802 21756 28812 21812
rect 28868 21756 28924 21812
rect 28980 21756 28990 21812
rect 31602 21756 31612 21812
rect 31668 21756 32172 21812
rect 32228 21756 33740 21812
rect 33796 21756 33806 21812
rect 34290 21756 34300 21812
rect 34356 21756 39340 21812
rect 39396 21756 39406 21812
rect 40450 21756 40460 21812
rect 40516 21756 41804 21812
rect 41860 21756 41870 21812
rect 27122 21644 27132 21700
rect 27188 21644 31276 21700
rect 31332 21644 31342 21700
rect 31714 21644 31724 21700
rect 31780 21644 33516 21700
rect 33572 21644 33582 21700
rect 38322 21644 38332 21700
rect 38388 21644 40236 21700
rect 40292 21644 40302 21700
rect 26338 21532 26348 21588
rect 26404 21532 26684 21588
rect 26740 21532 34076 21588
rect 34132 21532 34142 21588
rect 23426 21420 23436 21476
rect 23492 21420 24556 21476
rect 24612 21420 24622 21476
rect 25526 21420 25564 21476
rect 25620 21420 25630 21476
rect 28018 21420 28028 21476
rect 28084 21420 28094 21476
rect 30706 21420 30716 21476
rect 30772 21420 31724 21476
rect 31780 21420 31790 21476
rect 39330 21420 39340 21476
rect 39396 21420 41916 21476
rect 41972 21420 41982 21476
rect 22978 21308 22988 21364
rect 23044 21308 24108 21364
rect 24164 21308 25116 21364
rect 25172 21308 25182 21364
rect 28028 21252 28084 21420
rect 32610 21308 32620 21364
rect 32676 21308 33740 21364
rect 33796 21308 38444 21364
rect 38500 21308 38510 21364
rect 19618 21196 19628 21252
rect 19684 21196 28084 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 23426 21084 23436 21140
rect 23492 21084 34748 21140
rect 34804 21084 34814 21140
rect 27794 20972 27804 21028
rect 27860 20972 28140 21028
rect 28196 20972 38780 21028
rect 38836 20972 38846 21028
rect 1586 20860 1596 20916
rect 1652 20860 23884 20916
rect 23940 20860 23950 20916
rect 24332 20860 29596 20916
rect 29652 20860 29662 20916
rect 32722 20860 32732 20916
rect 32788 20860 33516 20916
rect 33572 20860 33582 20916
rect 34290 20860 34300 20916
rect 34356 20860 35756 20916
rect 35812 20860 36092 20916
rect 36148 20860 37996 20916
rect 38052 20860 38062 20916
rect 41570 20860 41580 20916
rect 41636 20860 42028 20916
rect 42084 20860 42364 20916
rect 42420 20860 42430 20916
rect 24332 20804 24388 20860
rect 22866 20748 22876 20804
rect 22932 20748 24388 20804
rect 26226 20748 26236 20804
rect 26292 20748 26684 20804
rect 26740 20748 36092 20804
rect 36148 20748 37436 20804
rect 37492 20748 37502 20804
rect 11330 20636 11340 20692
rect 11396 20636 24332 20692
rect 24388 20636 24398 20692
rect 26562 20636 26572 20692
rect 26628 20636 28700 20692
rect 28756 20636 29148 20692
rect 29204 20636 32732 20692
rect 32788 20636 32798 20692
rect 33506 20636 33516 20692
rect 33572 20636 36652 20692
rect 36708 20636 36718 20692
rect 21074 20524 21084 20580
rect 21140 20524 24668 20580
rect 24724 20524 27020 20580
rect 27076 20524 27086 20580
rect 27570 20524 27580 20580
rect 27636 20524 28588 20580
rect 28644 20524 29484 20580
rect 29540 20524 29550 20580
rect 30258 20524 30268 20580
rect 30324 20524 31836 20580
rect 31892 20524 31902 20580
rect 32610 20524 32620 20580
rect 32676 20524 33964 20580
rect 34020 20524 34300 20580
rect 34356 20524 34366 20580
rect 34738 20524 34748 20580
rect 34804 20524 35532 20580
rect 35588 20524 35598 20580
rect 35858 20524 35868 20580
rect 35924 20524 39228 20580
rect 39284 20524 39294 20580
rect 25778 20412 25788 20468
rect 25844 20412 27916 20468
rect 27972 20412 34916 20468
rect 36194 20412 36204 20468
rect 36260 20412 36540 20468
rect 36596 20412 40012 20468
rect 40068 20412 40078 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 34860 20356 34916 20412
rect 28354 20300 28364 20356
rect 28420 20300 28430 20356
rect 30706 20300 30716 20356
rect 30772 20300 33292 20356
rect 33348 20300 33358 20356
rect 34850 20300 34860 20356
rect 34916 20300 34926 20356
rect 36278 20300 36316 20356
rect 36372 20300 36382 20356
rect 36764 20300 39676 20356
rect 39732 20300 39742 20356
rect 20290 20188 20300 20244
rect 20356 20188 22876 20244
rect 22932 20188 22942 20244
rect 28364 20132 28420 20300
rect 36764 20244 36820 20300
rect 30594 20188 30604 20244
rect 30660 20188 31836 20244
rect 31892 20188 32620 20244
rect 32676 20188 32686 20244
rect 32834 20188 32844 20244
rect 32900 20188 36820 20244
rect 36978 20188 36988 20244
rect 37044 20188 37996 20244
rect 38052 20188 38062 20244
rect 25554 20076 25564 20132
rect 25620 20076 26124 20132
rect 26180 20076 27132 20132
rect 27188 20076 27198 20132
rect 28354 20076 28364 20132
rect 28420 20076 28430 20132
rect 33282 20076 33292 20132
rect 33348 20076 39340 20132
rect 39396 20076 39406 20132
rect 26002 19964 26012 20020
rect 26068 19964 27636 20020
rect 27794 19964 27804 20020
rect 27860 19964 28140 20020
rect 28196 19964 28206 20020
rect 28364 19964 33068 20020
rect 33124 19964 33134 20020
rect 33292 19964 33516 20020
rect 33572 19964 34412 20020
rect 34468 19964 34972 20020
rect 35028 19964 35038 20020
rect 37202 19964 37212 20020
rect 37268 19964 37884 20020
rect 37940 19964 37950 20020
rect 27580 19908 27636 19964
rect 28364 19908 28420 19964
rect 33292 19908 33348 19964
rect 22054 19852 22092 19908
rect 22148 19852 22158 19908
rect 24630 19852 24668 19908
rect 24724 19852 26124 19908
rect 26180 19852 27356 19908
rect 27412 19852 27422 19908
rect 27580 19852 28420 19908
rect 30146 19852 30156 19908
rect 30212 19852 31052 19908
rect 31108 19852 31118 19908
rect 32050 19852 32060 19908
rect 32116 19852 33348 19908
rect 33618 19852 33628 19908
rect 33684 19852 33964 19908
rect 34020 19852 34030 19908
rect 34962 19852 34972 19908
rect 35028 19852 35084 19908
rect 35140 19852 35150 19908
rect 36754 19852 36764 19908
rect 36820 19852 37100 19908
rect 37156 19852 37166 19908
rect 38406 19852 38444 19908
rect 38500 19852 38510 19908
rect 39106 19852 39116 19908
rect 39172 19852 40348 19908
rect 40404 19852 41468 19908
rect 41524 19852 41534 19908
rect 20962 19740 20972 19796
rect 21028 19740 24220 19796
rect 24276 19740 25900 19796
rect 25956 19740 25966 19796
rect 26898 19740 26908 19796
rect 26964 19740 27132 19796
rect 27188 19740 30044 19796
rect 30100 19740 30110 19796
rect 30818 19740 30828 19796
rect 30884 19740 30940 19796
rect 30996 19740 31388 19796
rect 31444 19740 31454 19796
rect 32610 19740 32620 19796
rect 32676 19740 36036 19796
rect 36194 19740 36204 19796
rect 36260 19740 36316 19796
rect 36372 19740 37996 19796
rect 38052 19740 40460 19796
rect 40516 19740 40526 19796
rect 35980 19684 36036 19740
rect 20738 19628 20748 19684
rect 20804 19628 27356 19684
rect 27412 19628 27422 19684
rect 27682 19628 27692 19684
rect 27748 19628 28252 19684
rect 28308 19628 28318 19684
rect 28578 19628 28588 19684
rect 28644 19628 29148 19684
rect 29204 19628 31948 19684
rect 32004 19628 32014 19684
rect 35980 19628 36988 19684
rect 37044 19628 37548 19684
rect 37604 19628 37614 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 22530 19516 22540 19572
rect 22596 19516 33012 19572
rect 35746 19516 35756 19572
rect 35812 19516 39788 19572
rect 39844 19516 39854 19572
rect 27122 19404 27132 19460
rect 27188 19404 28028 19460
rect 28084 19404 32284 19460
rect 32340 19404 32350 19460
rect 32956 19348 33012 19516
rect 33730 19404 33740 19460
rect 33796 19404 33852 19460
rect 33908 19404 41356 19460
rect 41412 19404 41422 19460
rect 28130 19292 28140 19348
rect 28196 19292 29148 19348
rect 29204 19292 29932 19348
rect 29988 19292 29998 19348
rect 32956 19292 34524 19348
rect 34580 19292 36764 19348
rect 36820 19292 36830 19348
rect 40674 19292 40684 19348
rect 40740 19292 42028 19348
rect 42084 19292 42094 19348
rect 41356 19236 41412 19292
rect 23650 19180 23660 19236
rect 23716 19180 25228 19236
rect 25284 19180 28028 19236
rect 28084 19180 28094 19236
rect 29586 19180 29596 19236
rect 29652 19180 32284 19236
rect 32340 19180 33516 19236
rect 33572 19180 33582 19236
rect 34178 19180 34188 19236
rect 34244 19180 34524 19236
rect 34580 19180 35532 19236
rect 35588 19180 35598 19236
rect 36390 19180 36428 19236
rect 36484 19180 36494 19236
rect 37538 19180 37548 19236
rect 37604 19180 38108 19236
rect 38164 19180 38174 19236
rect 41346 19180 41356 19236
rect 41412 19180 41422 19236
rect 24322 19068 24332 19124
rect 24388 19068 25004 19124
rect 25060 19068 25900 19124
rect 25956 19068 25966 19124
rect 27346 19068 27356 19124
rect 27412 19068 39676 19124
rect 39732 19068 39742 19124
rect 22194 18956 22204 19012
rect 22260 18956 22540 19012
rect 22596 18956 22606 19012
rect 25106 18956 25116 19012
rect 25172 18956 27132 19012
rect 27188 18956 27198 19012
rect 29362 18956 29372 19012
rect 29428 18956 29932 19012
rect 29988 18956 29998 19012
rect 31042 18956 31052 19012
rect 31108 18956 31500 19012
rect 31556 18956 31948 19012
rect 32834 18956 32844 19012
rect 32900 18956 33292 19012
rect 33348 18956 33358 19012
rect 35746 18956 35756 19012
rect 35812 18956 38108 19012
rect 38164 18956 39228 19012
rect 39284 18956 39294 19012
rect 40002 18956 40012 19012
rect 40068 18956 40684 19012
rect 40740 18956 40750 19012
rect 31892 18900 31948 18956
rect 30706 18844 30716 18900
rect 30772 18844 31612 18900
rect 31668 18844 31678 18900
rect 31892 18844 34524 18900
rect 34580 18844 34590 18900
rect 37398 18844 37436 18900
rect 37492 18844 37502 18900
rect 38770 18844 38780 18900
rect 38836 18844 38892 18900
rect 38948 18844 39900 18900
rect 39956 18844 39966 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 22978 18732 22988 18788
rect 23044 18732 27524 18788
rect 31938 18732 31948 18788
rect 32004 18732 35644 18788
rect 35700 18732 35710 18788
rect 27468 18676 27524 18732
rect 21634 18620 21644 18676
rect 21700 18620 24108 18676
rect 24164 18620 24174 18676
rect 26562 18620 26572 18676
rect 26628 18620 27132 18676
rect 27188 18620 27198 18676
rect 27468 18620 32620 18676
rect 32676 18620 32686 18676
rect 27132 18564 27188 18620
rect 18162 18508 18172 18564
rect 18228 18508 19852 18564
rect 19908 18508 23212 18564
rect 23268 18508 23278 18564
rect 23650 18508 23660 18564
rect 23716 18508 24332 18564
rect 24388 18508 24398 18564
rect 27132 18508 28140 18564
rect 28196 18508 28206 18564
rect 28466 18508 28476 18564
rect 28532 18508 28588 18564
rect 28644 18508 28654 18564
rect 30930 18508 30940 18564
rect 30996 18508 31164 18564
rect 31220 18508 31230 18564
rect 35830 18508 35868 18564
rect 35924 18508 35934 18564
rect 40450 18508 40460 18564
rect 40516 18508 40740 18564
rect 40684 18452 40740 18508
rect 20850 18396 20860 18452
rect 20916 18396 21532 18452
rect 21588 18396 21598 18452
rect 24210 18396 24220 18452
rect 24276 18396 26124 18452
rect 26180 18396 26684 18452
rect 26740 18396 27020 18452
rect 27076 18396 29484 18452
rect 29540 18396 29708 18452
rect 29764 18396 32396 18452
rect 32452 18396 32462 18452
rect 37762 18396 37772 18452
rect 37828 18396 39452 18452
rect 39508 18396 39518 18452
rect 40674 18396 40684 18452
rect 40740 18396 40750 18452
rect 1698 18284 1708 18340
rect 1764 18284 20076 18340
rect 20132 18284 20142 18340
rect 21298 18284 21308 18340
rect 21364 18284 21756 18340
rect 21812 18284 21822 18340
rect 30594 18284 30604 18340
rect 30660 18284 31052 18340
rect 31108 18284 31118 18340
rect 31602 18284 31612 18340
rect 31668 18284 32732 18340
rect 32788 18284 32798 18340
rect 32946 18284 32956 18340
rect 33012 18284 34076 18340
rect 34132 18284 34142 18340
rect 34850 18284 34860 18340
rect 34916 18284 35420 18340
rect 35476 18284 36652 18340
rect 36708 18284 36718 18340
rect 36866 18284 36876 18340
rect 36932 18284 37100 18340
rect 37156 18284 37660 18340
rect 37716 18284 37726 18340
rect 40786 18284 40796 18340
rect 40852 18284 41468 18340
rect 41524 18284 42028 18340
rect 42084 18284 42094 18340
rect 29250 18172 29260 18228
rect 29316 18172 30492 18228
rect 30548 18172 34132 18228
rect 34934 18172 34972 18228
rect 35028 18172 35980 18228
rect 36036 18172 36046 18228
rect 36418 18172 36428 18228
rect 36484 18172 39900 18228
rect 39956 18172 39966 18228
rect 41346 18172 41356 18228
rect 41412 18172 41804 18228
rect 41860 18172 41870 18228
rect 34076 18116 34132 18172
rect 28578 18060 28588 18116
rect 28644 18060 28924 18116
rect 28980 18060 29372 18116
rect 29428 18060 30044 18116
rect 30100 18060 31164 18116
rect 31220 18060 31948 18116
rect 32004 18060 32014 18116
rect 34066 18060 34076 18116
rect 34132 18060 34142 18116
rect 36642 18060 36652 18116
rect 36708 18060 38892 18116
rect 38948 18060 38958 18116
rect 41234 18060 41244 18116
rect 41300 18060 41916 18116
rect 41972 18060 41982 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 30492 18004 30548 18060
rect 31612 18004 31668 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19058 17948 19068 18004
rect 19124 17948 29820 18004
rect 29876 17948 30268 18004
rect 30324 17948 30334 18004
rect 30482 17948 30492 18004
rect 30548 17948 30558 18004
rect 31602 17948 31612 18004
rect 31668 17948 31678 18004
rect 37174 17948 37212 18004
rect 37268 17948 37278 18004
rect 41234 17948 41244 18004
rect 41300 17948 42364 18004
rect 42420 17948 42476 18004
rect 42532 17948 42542 18004
rect 25778 17836 25788 17892
rect 25844 17836 26236 17892
rect 26292 17836 27356 17892
rect 27412 17836 27422 17892
rect 34402 17836 34412 17892
rect 34468 17836 40460 17892
rect 40516 17836 40526 17892
rect 41356 17836 41692 17892
rect 41748 17836 41916 17892
rect 41972 17836 41982 17892
rect 41356 17780 41412 17836
rect 20850 17724 20860 17780
rect 20916 17724 21308 17780
rect 21364 17724 22092 17780
rect 22148 17724 22158 17780
rect 26002 17724 26012 17780
rect 26068 17724 30940 17780
rect 30996 17724 31006 17780
rect 31238 17724 31276 17780
rect 31332 17724 31342 17780
rect 40114 17724 40124 17780
rect 40180 17724 41412 17780
rect 41570 17724 41580 17780
rect 41636 17724 41916 17780
rect 41972 17724 41982 17780
rect 23762 17612 23772 17668
rect 23828 17612 24780 17668
rect 24836 17612 24846 17668
rect 30258 17612 30268 17668
rect 30324 17612 31500 17668
rect 31556 17612 31566 17668
rect 32498 17612 32508 17668
rect 32564 17612 33628 17668
rect 33684 17612 33694 17668
rect 38098 17612 38108 17668
rect 38164 17612 38388 17668
rect 24780 17556 24836 17612
rect 24780 17500 26572 17556
rect 26628 17500 26638 17556
rect 26898 17500 26908 17556
rect 26964 17500 27468 17556
rect 27524 17500 27534 17556
rect 31042 17500 31052 17556
rect 31108 17500 31556 17556
rect 31500 17444 31556 17500
rect 38332 17444 38388 17612
rect 38612 17612 42252 17668
rect 42308 17612 42318 17668
rect 26226 17388 26236 17444
rect 26292 17388 26684 17444
rect 26740 17388 26750 17444
rect 27346 17388 27356 17444
rect 27412 17388 28028 17444
rect 28084 17388 28094 17444
rect 30146 17388 30156 17444
rect 30212 17388 31276 17444
rect 31332 17388 31342 17444
rect 31490 17388 31500 17444
rect 31556 17388 31566 17444
rect 33058 17388 33068 17444
rect 33124 17388 38108 17444
rect 38164 17388 38174 17444
rect 38322 17388 38332 17444
rect 38388 17388 38444 17444
rect 38500 17388 38510 17444
rect 38612 17332 38668 17612
rect 38994 17388 39004 17444
rect 39060 17388 39340 17444
rect 39396 17388 39406 17444
rect 41318 17388 41356 17444
rect 41412 17388 41422 17444
rect 21756 17276 25564 17332
rect 25620 17276 25630 17332
rect 27234 17276 27244 17332
rect 27300 17276 31948 17332
rect 33954 17276 33964 17332
rect 34020 17276 34636 17332
rect 34692 17276 38668 17332
rect 40450 17276 40460 17332
rect 40516 17276 41916 17332
rect 41972 17276 41982 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 17266 17164 17276 17220
rect 17332 17164 19516 17220
rect 19572 17164 19582 17220
rect 20178 17164 20188 17220
rect 20244 17164 21084 17220
rect 21140 17164 21150 17220
rect 21756 17108 21812 17276
rect 21970 17164 21980 17220
rect 22036 17164 25564 17220
rect 25620 17164 25630 17220
rect 29810 17164 29820 17220
rect 29876 17164 30604 17220
rect 30660 17164 31724 17220
rect 31780 17164 31790 17220
rect 18722 17052 18732 17108
rect 18788 17052 21812 17108
rect 23986 17052 23996 17108
rect 24052 17052 24062 17108
rect 17612 16940 18788 16996
rect 19506 16940 19516 16996
rect 19572 16940 21308 16996
rect 21364 16940 21374 16996
rect 21746 16940 21756 16996
rect 21812 16940 22988 16996
rect 23044 16940 23054 16996
rect 17612 16884 17668 16940
rect 18732 16884 18788 16940
rect 23996 16884 24052 17052
rect 26450 16940 26460 16996
rect 26516 16940 27244 16996
rect 27300 16940 27310 16996
rect 27570 16940 27580 16996
rect 27636 16940 28476 16996
rect 28532 16940 28542 16996
rect 15250 16828 15260 16884
rect 15316 16828 15484 16884
rect 15540 16828 15550 16884
rect 16930 16828 16940 16884
rect 16996 16828 17612 16884
rect 17668 16828 17678 16884
rect 18274 16828 18284 16884
rect 18340 16828 18508 16884
rect 18564 16828 18574 16884
rect 18732 16828 24052 16884
rect 25554 16828 25564 16884
rect 25620 16828 26348 16884
rect 26404 16828 26414 16884
rect 26562 16828 26572 16884
rect 26628 16828 27020 16884
rect 27076 16828 27086 16884
rect 28354 16828 28364 16884
rect 28420 16828 29036 16884
rect 29092 16828 29102 16884
rect 29820 16772 29876 17164
rect 31892 17108 31948 17276
rect 32050 17164 32060 17220
rect 32116 17164 32620 17220
rect 32676 17164 32686 17220
rect 33618 17164 33628 17220
rect 33684 17164 34748 17220
rect 34804 17164 40012 17220
rect 40068 17164 40572 17220
rect 40628 17164 41580 17220
rect 41636 17164 41646 17220
rect 31892 17052 32172 17108
rect 32228 17052 36204 17108
rect 36260 17052 36270 17108
rect 36530 17052 36540 17108
rect 36596 17052 37100 17108
rect 37156 17052 37166 17108
rect 37314 17052 37324 17108
rect 37380 17052 38668 17108
rect 38724 17052 38734 17108
rect 41206 17052 41244 17108
rect 41300 17052 41310 17108
rect 30370 16940 30380 16996
rect 30436 16940 31388 16996
rect 31444 16940 31454 16996
rect 32386 16940 32396 16996
rect 32452 16940 33740 16996
rect 33796 16940 33806 16996
rect 36306 16940 36316 16996
rect 36372 16940 38332 16996
rect 38388 16940 39116 16996
rect 39172 16940 39788 16996
rect 39844 16940 40572 16996
rect 40628 16940 40638 16996
rect 43138 16940 43148 16996
rect 43204 16940 43214 16996
rect 43148 16884 43204 16940
rect 32722 16828 32732 16884
rect 32788 16828 34412 16884
rect 34468 16828 34478 16884
rect 36642 16828 36652 16884
rect 36708 16828 37324 16884
rect 37380 16828 37390 16884
rect 37986 16828 37996 16884
rect 38052 16828 39340 16884
rect 39396 16828 39406 16884
rect 39666 16828 39676 16884
rect 39732 16828 40460 16884
rect 40516 16828 40526 16884
rect 41804 16828 43372 16884
rect 43428 16828 43438 16884
rect 41804 16772 41860 16828
rect 19058 16716 19068 16772
rect 19124 16716 22428 16772
rect 22484 16716 22494 16772
rect 22642 16716 22652 16772
rect 22708 16716 23324 16772
rect 23380 16716 28476 16772
rect 28532 16716 28542 16772
rect 28914 16716 28924 16772
rect 28980 16716 29932 16772
rect 29988 16716 29998 16772
rect 41794 16716 41804 16772
rect 41860 16716 41870 16772
rect 22652 16660 22708 16716
rect 20178 16604 20188 16660
rect 20244 16604 22708 16660
rect 24882 16604 24892 16660
rect 24948 16604 25900 16660
rect 25956 16604 25966 16660
rect 31266 16604 31276 16660
rect 31332 16604 31724 16660
rect 31780 16604 32844 16660
rect 32900 16604 35588 16660
rect 39218 16604 39228 16660
rect 39284 16604 41020 16660
rect 41076 16604 41692 16660
rect 41748 16604 41758 16660
rect 35532 16548 35588 16604
rect 27458 16492 27468 16548
rect 27524 16492 28364 16548
rect 28420 16492 28430 16548
rect 29586 16492 29596 16548
rect 29652 16492 30044 16548
rect 30100 16492 30716 16548
rect 30772 16492 30782 16548
rect 33254 16492 33292 16548
rect 33348 16492 33358 16548
rect 35532 16492 40348 16548
rect 40404 16492 40414 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 27346 16380 27356 16436
rect 27412 16380 27804 16436
rect 27860 16380 27870 16436
rect 28214 16380 28252 16436
rect 28308 16380 28318 16436
rect 31826 16380 31836 16436
rect 31892 16380 33852 16436
rect 33908 16380 33918 16436
rect 35634 16380 35644 16436
rect 35700 16380 35980 16436
rect 36036 16380 36046 16436
rect 36194 16380 36204 16436
rect 36260 16380 36764 16436
rect 36820 16380 36830 16436
rect 38658 16380 38668 16436
rect 38724 16380 39900 16436
rect 39956 16380 39966 16436
rect 41878 16380 41916 16436
rect 41972 16380 41982 16436
rect 18722 16268 18732 16324
rect 18788 16268 20412 16324
rect 20468 16268 20478 16324
rect 24210 16268 24220 16324
rect 24276 16268 24286 16324
rect 25106 16268 25116 16324
rect 25172 16268 41468 16324
rect 41524 16268 41534 16324
rect 24220 16212 24276 16268
rect 19170 16156 19180 16212
rect 19236 16156 20860 16212
rect 20916 16156 20926 16212
rect 22306 16156 22316 16212
rect 22372 16156 23212 16212
rect 23268 16156 23278 16212
rect 24220 16156 24668 16212
rect 24724 16156 26348 16212
rect 26404 16156 31164 16212
rect 31220 16156 31230 16212
rect 33394 16156 33404 16212
rect 33460 16156 33628 16212
rect 33684 16156 33694 16212
rect 34962 16156 34972 16212
rect 35028 16156 35308 16212
rect 35364 16156 35756 16212
rect 35812 16156 36540 16212
rect 36596 16156 36606 16212
rect 37426 16156 37436 16212
rect 37492 16156 39564 16212
rect 39620 16156 39630 16212
rect 23100 16044 23436 16100
rect 23492 16044 24108 16100
rect 24164 16044 24174 16100
rect 24322 16044 24332 16100
rect 24388 16044 24780 16100
rect 24836 16044 25452 16100
rect 25508 16044 25518 16100
rect 25890 16044 25900 16100
rect 25956 16044 28252 16100
rect 28308 16044 28588 16100
rect 28644 16044 28654 16100
rect 30930 16044 30940 16100
rect 30996 16044 31836 16100
rect 31892 16044 31902 16100
rect 32498 16044 32508 16100
rect 32564 16044 32844 16100
rect 32900 16044 32910 16100
rect 36306 16044 36316 16100
rect 36372 16044 37660 16100
rect 37716 16044 37726 16100
rect 39078 16044 39116 16100
rect 39172 16044 39182 16100
rect 39330 16044 39340 16100
rect 39396 16044 41468 16100
rect 41524 16044 41804 16100
rect 41860 16044 41870 16100
rect 23100 15988 23156 16044
rect 23090 15932 23100 15988
rect 23156 15932 23166 15988
rect 27318 15932 27356 15988
rect 27412 15932 27422 15988
rect 28242 15932 28252 15988
rect 28308 15932 28364 15988
rect 28420 15932 28430 15988
rect 31490 15932 31500 15988
rect 31556 15932 32956 15988
rect 33012 15932 33022 15988
rect 34738 15932 34748 15988
rect 34804 15932 34860 15988
rect 34916 15932 35420 15988
rect 35476 15932 35486 15988
rect 36530 15932 36540 15988
rect 36596 15932 37212 15988
rect 37268 15932 37278 15988
rect 38882 15932 38892 15988
rect 38948 15932 39452 15988
rect 39508 15932 39518 15988
rect 40534 15932 40572 15988
rect 40628 15932 40638 15988
rect 6738 15820 6748 15876
rect 6804 15820 15708 15876
rect 15764 15820 15774 15876
rect 16034 15820 16044 15876
rect 16100 15820 17948 15876
rect 18004 15820 21644 15876
rect 21700 15820 22204 15876
rect 22260 15820 22270 15876
rect 23426 15820 23436 15876
rect 23492 15820 24220 15876
rect 24276 15820 24286 15876
rect 29810 15820 29820 15876
rect 29876 15820 30044 15876
rect 30100 15820 30110 15876
rect 34402 15820 34412 15876
rect 34468 15820 36316 15876
rect 36372 15820 36382 15876
rect 36642 15820 36652 15876
rect 36708 15820 38052 15876
rect 39890 15820 39900 15876
rect 39956 15820 41020 15876
rect 41076 15820 41086 15876
rect 41458 15820 41468 15876
rect 41524 15820 41692 15876
rect 41748 15820 41758 15876
rect 22204 15764 22260 15820
rect 37996 15764 38052 15820
rect 22204 15708 26236 15764
rect 26292 15708 27020 15764
rect 27076 15708 27086 15764
rect 28466 15708 28476 15764
rect 28532 15708 29764 15764
rect 30146 15708 30156 15764
rect 30212 15708 35476 15764
rect 35634 15708 35644 15764
rect 35700 15708 37212 15764
rect 37268 15708 37772 15764
rect 37828 15708 37838 15764
rect 37996 15708 40012 15764
rect 40068 15708 40078 15764
rect 40338 15708 40348 15764
rect 40404 15708 40572 15764
rect 40628 15708 40638 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 29708 15652 29764 15708
rect 35420 15652 35476 15708
rect 26898 15596 26908 15652
rect 26964 15596 29484 15652
rect 29540 15596 29550 15652
rect 29708 15596 32172 15652
rect 32228 15596 32284 15652
rect 32340 15596 32620 15652
rect 32676 15596 32686 15652
rect 32834 15596 32844 15652
rect 32900 15596 32910 15652
rect 35420 15596 35924 15652
rect 36642 15596 36652 15652
rect 36708 15596 37436 15652
rect 37492 15596 37502 15652
rect 38210 15596 38220 15652
rect 38276 15596 40460 15652
rect 40516 15596 40526 15652
rect 32844 15540 32900 15596
rect 35868 15540 35924 15596
rect 13346 15484 13356 15540
rect 13412 15484 14364 15540
rect 14420 15484 14430 15540
rect 15698 15484 15708 15540
rect 15764 15484 19964 15540
rect 20020 15484 20030 15540
rect 27122 15484 27132 15540
rect 27188 15484 28140 15540
rect 28196 15484 28206 15540
rect 29586 15484 29596 15540
rect 29652 15484 30380 15540
rect 30436 15484 30446 15540
rect 30594 15484 30604 15540
rect 30660 15484 31388 15540
rect 31444 15484 31454 15540
rect 32844 15484 34636 15540
rect 34692 15484 35644 15540
rect 35700 15484 35710 15540
rect 35868 15484 36764 15540
rect 36820 15484 36830 15540
rect 39442 15484 39452 15540
rect 39508 15484 40236 15540
rect 40292 15484 40302 15540
rect 30604 15428 30660 15484
rect 21298 15372 21308 15428
rect 21364 15372 21980 15428
rect 22036 15372 22046 15428
rect 22418 15372 22428 15428
rect 22484 15372 23324 15428
rect 23380 15372 24668 15428
rect 24724 15372 25116 15428
rect 25172 15372 25676 15428
rect 25732 15372 28588 15428
rect 28644 15372 28654 15428
rect 29474 15372 29484 15428
rect 29540 15372 30660 15428
rect 32162 15372 32172 15428
rect 32228 15372 34916 15428
rect 36306 15372 36316 15428
rect 36372 15372 37100 15428
rect 37156 15372 37166 15428
rect 37426 15372 37436 15428
rect 37492 15372 38332 15428
rect 38388 15372 38398 15428
rect 38546 15372 38556 15428
rect 38612 15372 39564 15428
rect 39620 15372 39630 15428
rect 34860 15316 34916 15372
rect 26002 15260 26012 15316
rect 26068 15260 26796 15316
rect 26852 15260 26862 15316
rect 27458 15260 27468 15316
rect 27524 15260 29372 15316
rect 29428 15260 29438 15316
rect 29698 15260 29708 15316
rect 29764 15260 30268 15316
rect 30324 15260 30716 15316
rect 30772 15260 32284 15316
rect 32340 15260 32350 15316
rect 32498 15260 32508 15316
rect 32564 15260 33516 15316
rect 33572 15260 33582 15316
rect 33730 15260 33740 15316
rect 33796 15260 34076 15316
rect 34132 15260 34142 15316
rect 34850 15260 34860 15316
rect 34916 15260 35532 15316
rect 35588 15260 35598 15316
rect 36418 15260 36428 15316
rect 36484 15260 38444 15316
rect 38500 15260 38510 15316
rect 38770 15260 38780 15316
rect 38836 15260 40236 15316
rect 40292 15260 40302 15316
rect 40674 15260 40684 15316
rect 40740 15260 41692 15316
rect 41748 15260 41758 15316
rect 10098 15148 10108 15204
rect 10164 15148 12572 15204
rect 12628 15148 13916 15204
rect 13972 15148 15820 15204
rect 15876 15148 15886 15204
rect 27234 15148 27244 15204
rect 27300 15148 28812 15204
rect 28868 15148 28878 15204
rect 29036 15148 29484 15204
rect 29540 15148 29550 15204
rect 31490 15148 31500 15204
rect 31556 15148 32396 15204
rect 32452 15148 33964 15204
rect 34020 15148 34030 15204
rect 35634 15148 35644 15204
rect 35700 15148 35868 15204
rect 35924 15148 35934 15204
rect 41458 15148 41468 15204
rect 41524 15148 41804 15204
rect 41860 15148 41870 15204
rect 29036 15092 29092 15148
rect 9650 15036 9660 15092
rect 9716 15036 17500 15092
rect 17556 15036 17566 15092
rect 22978 15036 22988 15092
rect 23044 15036 23548 15092
rect 23604 15036 25228 15092
rect 25284 15036 27020 15092
rect 27076 15036 28028 15092
rect 28084 15036 28094 15092
rect 28466 15036 28476 15092
rect 28532 15036 29092 15092
rect 8418 14924 8428 14980
rect 8484 14924 18620 14980
rect 18676 14924 20076 14980
rect 20132 14924 20142 14980
rect 32134 14924 32172 14980
rect 32228 14924 32238 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 16594 14812 16604 14868
rect 16660 14812 25564 14868
rect 25620 14812 26348 14868
rect 26404 14812 26414 14868
rect 28438 14812 28476 14868
rect 28532 14812 28542 14868
rect 30818 14812 30828 14868
rect 30884 14812 34860 14868
rect 34916 14812 34926 14868
rect 38658 14812 38668 14868
rect 38724 14812 38892 14868
rect 38948 14812 38958 14868
rect 28690 14700 28700 14756
rect 28756 14700 31276 14756
rect 31332 14700 31342 14756
rect 33506 14700 33516 14756
rect 33572 14700 33852 14756
rect 33908 14700 33918 14756
rect 16482 14588 16492 14644
rect 16548 14588 18172 14644
rect 18228 14588 18238 14644
rect 28028 14588 29036 14644
rect 29092 14588 29102 14644
rect 31378 14588 31388 14644
rect 31444 14588 33292 14644
rect 33348 14588 33358 14644
rect 33618 14588 33628 14644
rect 33684 14588 37100 14644
rect 37156 14588 37324 14644
rect 37380 14588 37390 14644
rect 39890 14588 39900 14644
rect 39956 14588 40236 14644
rect 40292 14588 40302 14644
rect 17938 14476 17948 14532
rect 18004 14476 19628 14532
rect 19684 14476 19694 14532
rect 25890 14476 25900 14532
rect 25956 14476 26572 14532
rect 26628 14476 26638 14532
rect 27094 14476 27132 14532
rect 27188 14476 27198 14532
rect 15474 14364 15484 14420
rect 15540 14364 19516 14420
rect 19572 14364 21420 14420
rect 21476 14364 21486 14420
rect 25218 14364 25228 14420
rect 25284 14364 27300 14420
rect 27244 14308 27300 14364
rect 28028 14308 28084 14588
rect 28578 14476 28588 14532
rect 28644 14476 29148 14532
rect 29204 14476 29214 14532
rect 29698 14476 29708 14532
rect 29764 14476 30492 14532
rect 30548 14476 30558 14532
rect 32610 14476 32620 14532
rect 32676 14476 36204 14532
rect 36260 14476 36270 14532
rect 41878 14476 41916 14532
rect 41972 14476 41982 14532
rect 28802 14364 28812 14420
rect 28868 14364 30604 14420
rect 30660 14364 32060 14420
rect 32116 14364 34300 14420
rect 34356 14364 34524 14420
rect 34580 14364 34590 14420
rect 39106 14364 39116 14420
rect 39172 14364 39564 14420
rect 39620 14364 39630 14420
rect 39890 14364 39900 14420
rect 39956 14364 40684 14420
rect 40740 14364 40750 14420
rect 15250 14252 15260 14308
rect 15316 14252 15596 14308
rect 15652 14252 15662 14308
rect 17042 14252 17052 14308
rect 17108 14252 17388 14308
rect 17444 14252 17454 14308
rect 18834 14252 18844 14308
rect 18900 14252 20244 14308
rect 20850 14252 20860 14308
rect 20916 14252 21756 14308
rect 21812 14252 24220 14308
rect 24276 14252 25900 14308
rect 25956 14252 25966 14308
rect 27234 14252 27244 14308
rect 27300 14252 28028 14308
rect 28084 14252 28094 14308
rect 28914 14252 28924 14308
rect 28980 14252 30492 14308
rect 30548 14252 30558 14308
rect 31948 14252 36652 14308
rect 36708 14252 37436 14308
rect 37492 14252 38108 14308
rect 38164 14252 38174 14308
rect 41346 14252 41356 14308
rect 41412 14252 41692 14308
rect 41748 14252 41758 14308
rect 20188 14196 20244 14252
rect 15138 14140 15148 14196
rect 15204 14140 17164 14196
rect 17220 14140 17230 14196
rect 20178 14140 20188 14196
rect 20244 14140 20254 14196
rect 29026 14140 29036 14196
rect 29092 14140 31388 14196
rect 31444 14140 31454 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 31948 14084 32004 14252
rect 33842 14140 33852 14196
rect 33908 14140 34972 14196
rect 35028 14140 38444 14196
rect 38500 14140 38510 14196
rect 40674 14140 40684 14196
rect 40740 14140 41580 14196
rect 41636 14140 41646 14196
rect 14252 14028 19068 14084
rect 19124 14028 19134 14084
rect 20402 14028 20412 14084
rect 20468 14028 21644 14084
rect 21700 14028 21710 14084
rect 28578 14028 28588 14084
rect 28644 14028 29596 14084
rect 29652 14028 32004 14084
rect 32162 14028 32172 14084
rect 32228 14028 33628 14084
rect 33684 14028 37772 14084
rect 37828 14028 37838 14084
rect 42326 14028 42364 14084
rect 42420 14028 42430 14084
rect 14252 13860 14308 14028
rect 16828 13916 16940 13972
rect 16996 13916 17948 13972
rect 18004 13916 18014 13972
rect 6402 13804 6412 13860
rect 6468 13804 9100 13860
rect 9156 13804 11116 13860
rect 11172 13804 11182 13860
rect 12898 13804 12908 13860
rect 12964 13804 13132 13860
rect 13188 13804 14252 13860
rect 14308 13804 14318 13860
rect 14914 13804 14924 13860
rect 14980 13804 15148 13860
rect 15204 13804 15214 13860
rect 16828 13748 16884 13916
rect 19068 13860 19124 14028
rect 19618 13916 19628 13972
rect 19684 13916 25452 13972
rect 25508 13916 25518 13972
rect 27234 13916 27244 13972
rect 27300 13916 28364 13972
rect 28420 13916 32564 13972
rect 32834 13916 32844 13972
rect 32900 13916 33852 13972
rect 33908 13916 37548 13972
rect 37604 13916 37614 13972
rect 39488 13916 39564 13972
rect 39620 13916 40572 13972
rect 40628 13916 40638 13972
rect 41654 13916 41692 13972
rect 41748 13916 41758 13972
rect 21532 13860 21588 13916
rect 32508 13860 32564 13916
rect 19068 13804 21308 13860
rect 21364 13804 21374 13860
rect 21522 13804 21532 13860
rect 21588 13804 21598 13860
rect 23202 13804 23212 13860
rect 23268 13804 28476 13860
rect 28532 13804 28542 13860
rect 29922 13804 29932 13860
rect 29988 13804 30492 13860
rect 30548 13804 30558 13860
rect 32498 13804 32508 13860
rect 32564 13804 35812 13860
rect 35970 13804 35980 13860
rect 36036 13804 37212 13860
rect 37268 13804 37772 13860
rect 37828 13804 37838 13860
rect 38322 13804 38332 13860
rect 38388 13804 39676 13860
rect 39732 13804 39742 13860
rect 25900 13748 25956 13804
rect 35756 13748 35812 13804
rect 3938 13692 3948 13748
rect 4004 13692 13356 13748
rect 13412 13692 13692 13748
rect 13748 13692 13758 13748
rect 14690 13692 14700 13748
rect 14756 13692 16884 13748
rect 17378 13692 17388 13748
rect 17444 13692 17836 13748
rect 17892 13692 19180 13748
rect 19236 13692 19740 13748
rect 19796 13692 19806 13748
rect 20402 13692 20412 13748
rect 20468 13692 20972 13748
rect 21028 13692 23492 13748
rect 24434 13692 24444 13748
rect 24500 13692 24780 13748
rect 24836 13692 24846 13748
rect 25442 13692 25452 13748
rect 25508 13692 25676 13748
rect 25732 13692 25742 13748
rect 25890 13692 25900 13748
rect 25956 13692 25966 13748
rect 26338 13692 26348 13748
rect 26404 13692 26908 13748
rect 26964 13692 26974 13748
rect 27346 13692 27356 13748
rect 27412 13692 30492 13748
rect 30548 13692 32732 13748
rect 32788 13692 32798 13748
rect 33254 13692 33292 13748
rect 33348 13692 33358 13748
rect 34290 13692 34300 13748
rect 34356 13692 35532 13748
rect 35588 13692 35598 13748
rect 35756 13692 36540 13748
rect 36596 13692 36764 13748
rect 36820 13692 36830 13748
rect 38182 13692 38220 13748
rect 38276 13692 38286 13748
rect 40562 13692 40572 13748
rect 40628 13692 41244 13748
rect 41300 13692 42588 13748
rect 42644 13692 42654 13748
rect 13692 13636 13748 13692
rect 23436 13636 23492 13692
rect 2930 13580 2940 13636
rect 2996 13580 3388 13636
rect 8978 13580 8988 13636
rect 9044 13580 10332 13636
rect 10388 13580 10398 13636
rect 12002 13580 12012 13636
rect 12068 13580 12908 13636
rect 12964 13580 12974 13636
rect 13692 13580 14924 13636
rect 14980 13580 14990 13636
rect 15698 13580 15708 13636
rect 15764 13580 16044 13636
rect 16100 13580 17612 13636
rect 17668 13580 17678 13636
rect 18610 13580 18620 13636
rect 18676 13580 22764 13636
rect 22820 13580 22830 13636
rect 23426 13580 23436 13636
rect 23492 13580 24388 13636
rect 24546 13580 24556 13636
rect 24612 13580 25788 13636
rect 25844 13580 25854 13636
rect 3332 13524 3388 13580
rect 24332 13524 24388 13580
rect 27356 13524 27412 13692
rect 28018 13580 28028 13636
rect 28084 13580 29372 13636
rect 29428 13580 29438 13636
rect 32050 13580 32060 13636
rect 32116 13580 33628 13636
rect 33684 13580 33694 13636
rect 34738 13580 34748 13636
rect 34804 13580 34972 13636
rect 35028 13580 35038 13636
rect 38098 13580 38108 13636
rect 38164 13580 40684 13636
rect 40740 13580 40750 13636
rect 3332 13468 13916 13524
rect 13972 13468 13982 13524
rect 18386 13468 18396 13524
rect 18452 13468 23660 13524
rect 23716 13468 23726 13524
rect 24332 13468 27412 13524
rect 29250 13468 29260 13524
rect 29316 13468 29820 13524
rect 29876 13468 32396 13524
rect 32452 13468 35420 13524
rect 35476 13468 35486 13524
rect 35858 13468 35868 13524
rect 35924 13468 36652 13524
rect 36708 13468 36988 13524
rect 37044 13468 38108 13524
rect 38164 13468 38174 13524
rect 22642 13356 22652 13412
rect 22708 13356 23548 13412
rect 23604 13356 23614 13412
rect 24630 13356 24668 13412
rect 24724 13356 24734 13412
rect 24882 13356 24892 13412
rect 24948 13356 28364 13412
rect 28420 13356 28588 13412
rect 28644 13356 28654 13412
rect 30818 13356 30828 13412
rect 30884 13356 32284 13412
rect 32340 13356 32350 13412
rect 33058 13356 33068 13412
rect 33124 13356 33964 13412
rect 34020 13356 34030 13412
rect 34850 13356 34860 13412
rect 34916 13356 34972 13412
rect 35028 13356 35038 13412
rect 39330 13356 39340 13412
rect 39396 13356 40012 13412
rect 40068 13356 40572 13412
rect 40628 13356 40638 13412
rect 41570 13356 41580 13412
rect 41636 13356 41916 13412
rect 41972 13356 41982 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 5954 13244 5964 13300
rect 6020 13244 7196 13300
rect 7252 13244 14588 13300
rect 14644 13244 14654 13300
rect 15092 13244 20636 13300
rect 20692 13244 21084 13300
rect 21140 13244 21150 13300
rect 26226 13244 26236 13300
rect 26292 13244 28252 13300
rect 28308 13244 28318 13300
rect 29138 13244 29148 13300
rect 29204 13244 33852 13300
rect 33908 13244 33918 13300
rect 36306 13244 36316 13300
rect 36372 13244 37324 13300
rect 37380 13244 37390 13300
rect 41682 13244 41692 13300
rect 41748 13244 42140 13300
rect 42196 13244 42206 13300
rect 15092 13076 15148 13244
rect 19394 13132 19404 13188
rect 19460 13132 22316 13188
rect 22372 13132 22382 13188
rect 28466 13132 28476 13188
rect 28532 13132 38780 13188
rect 38836 13132 40012 13188
rect 40068 13132 40078 13188
rect 3332 13020 15148 13076
rect 21970 13020 21980 13076
rect 22036 13020 22988 13076
rect 23044 13020 23054 13076
rect 26002 13020 26012 13076
rect 26068 13020 26796 13076
rect 26852 13020 27132 13076
rect 27188 13020 27198 13076
rect 27346 13020 27356 13076
rect 27412 13020 30828 13076
rect 30884 13020 30894 13076
rect 31042 13020 31052 13076
rect 31108 13020 32060 13076
rect 32116 13020 33516 13076
rect 33572 13020 33582 13076
rect 33954 13020 33964 13076
rect 34020 13020 35196 13076
rect 35252 13020 35756 13076
rect 35812 13020 37660 13076
rect 37716 13020 39116 13076
rect 39172 13020 39182 13076
rect 42242 13020 42252 13076
rect 42308 13020 42812 13076
rect 42868 13020 42878 13076
rect 3332 12628 3388 13020
rect 14578 12908 14588 12964
rect 14644 12908 15036 12964
rect 15092 12908 15102 12964
rect 28690 12908 28700 12964
rect 28756 12908 30156 12964
rect 30212 12908 30222 12964
rect 30370 12908 30380 12964
rect 30436 12908 31892 12964
rect 32834 12908 32844 12964
rect 32900 12908 36988 12964
rect 37044 12908 37054 12964
rect 38546 12908 38556 12964
rect 38612 12908 38668 12964
rect 38724 12908 38734 12964
rect 39666 12908 39676 12964
rect 39732 12908 40572 12964
rect 40628 12908 40638 12964
rect 41430 12908 41468 12964
rect 41524 12908 41534 12964
rect 31836 12852 31892 12908
rect 11218 12796 11228 12852
rect 11284 12796 12012 12852
rect 12068 12796 12078 12852
rect 17266 12796 17276 12852
rect 17332 12796 21980 12852
rect 22036 12796 22988 12852
rect 23044 12796 24892 12852
rect 24948 12796 24958 12852
rect 26562 12796 26572 12852
rect 26628 12796 27692 12852
rect 27748 12796 27758 12852
rect 28354 12796 28364 12852
rect 28420 12796 30604 12852
rect 30660 12796 30670 12852
rect 31574 12796 31612 12852
rect 31668 12796 31678 12852
rect 31836 12796 34300 12852
rect 34356 12796 34366 12852
rect 36082 12796 36092 12852
rect 36148 12796 36764 12852
rect 36820 12796 37324 12852
rect 37380 12796 37390 12852
rect 37650 12796 37660 12852
rect 37716 12796 38108 12852
rect 38164 12796 39004 12852
rect 39060 12796 39900 12852
rect 39956 12796 39966 12852
rect 8530 12684 8540 12740
rect 8596 12684 10668 12740
rect 10724 12684 10734 12740
rect 11442 12684 11452 12740
rect 11508 12684 12796 12740
rect 12852 12684 12862 12740
rect 13468 12684 13804 12740
rect 13860 12684 13870 12740
rect 14354 12684 14364 12740
rect 14420 12684 16268 12740
rect 16324 12684 18844 12740
rect 18900 12684 18910 12740
rect 24322 12684 24332 12740
rect 24388 12684 25900 12740
rect 25956 12684 28140 12740
rect 28196 12684 28206 12740
rect 30706 12684 30716 12740
rect 30772 12684 30940 12740
rect 30996 12684 31006 12740
rect 31490 12684 31500 12740
rect 31556 12684 33740 12740
rect 33796 12684 34748 12740
rect 34804 12684 34814 12740
rect 37762 12684 37772 12740
rect 37828 12684 38780 12740
rect 38836 12684 38846 12740
rect 39778 12684 39788 12740
rect 39844 12684 40684 12740
rect 40740 12684 42028 12740
rect 42084 12684 42094 12740
rect 13468 12628 13524 12684
rect 2034 12572 2044 12628
rect 2100 12572 3388 12628
rect 12338 12572 12348 12628
rect 12404 12572 12908 12628
rect 12964 12572 13468 12628
rect 13524 12572 13534 12628
rect 13682 12572 13692 12628
rect 13748 12572 13916 12628
rect 13972 12572 14476 12628
rect 14532 12572 14542 12628
rect 14802 12572 14812 12628
rect 14868 12572 14878 12628
rect 15474 12572 15484 12628
rect 15540 12572 18732 12628
rect 18788 12572 18798 12628
rect 26674 12572 26684 12628
rect 26740 12572 26908 12628
rect 26964 12572 26974 12628
rect 29922 12572 29932 12628
rect 29988 12572 31948 12628
rect 32004 12572 32014 12628
rect 36194 12572 36204 12628
rect 36260 12572 40572 12628
rect 40628 12572 40638 12628
rect 41682 12572 41692 12628
rect 41748 12572 41758 12628
rect 14812 12516 14868 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 31948 12516 32004 12572
rect 41692 12516 41748 12572
rect 9874 12460 9884 12516
rect 9940 12460 9950 12516
rect 11554 12460 11564 12516
rect 11620 12460 12460 12516
rect 12516 12460 12526 12516
rect 14476 12460 14868 12516
rect 30678 12460 30716 12516
rect 30772 12460 30782 12516
rect 30930 12460 30940 12516
rect 30996 12460 31052 12516
rect 31108 12460 31118 12516
rect 31948 12460 36428 12516
rect 36484 12460 36494 12516
rect 37202 12460 37212 12516
rect 37268 12460 41748 12516
rect 9884 12404 9940 12460
rect 9426 12348 9436 12404
rect 9492 12348 10220 12404
rect 10276 12348 10286 12404
rect 11106 12348 11116 12404
rect 11172 12348 12796 12404
rect 12852 12348 12862 12404
rect 9314 12236 9324 12292
rect 9380 12236 9884 12292
rect 9940 12236 9950 12292
rect 10322 12236 10332 12292
rect 10388 12236 14252 12292
rect 14308 12236 14318 12292
rect 10332 12180 10388 12236
rect 14476 12180 14532 12460
rect 14802 12348 14812 12404
rect 14868 12348 15148 12404
rect 15204 12348 15214 12404
rect 15810 12348 15820 12404
rect 15876 12348 18676 12404
rect 29782 12348 29820 12404
rect 29876 12348 31388 12404
rect 31444 12348 31454 12404
rect 31602 12348 31612 12404
rect 31668 12348 33516 12404
rect 33572 12348 36652 12404
rect 36708 12348 36718 12404
rect 38322 12348 38332 12404
rect 38388 12348 38444 12404
rect 38500 12348 38510 12404
rect 39442 12348 39452 12404
rect 39508 12348 39564 12404
rect 39620 12348 39630 12404
rect 41010 12348 41020 12404
rect 41076 12348 41692 12404
rect 41748 12348 41758 12404
rect 16818 12236 16828 12292
rect 16884 12236 17052 12292
rect 17108 12236 17118 12292
rect 18620 12180 18676 12348
rect 18834 12236 18844 12292
rect 18900 12236 20412 12292
rect 20468 12236 20478 12292
rect 27542 12236 27580 12292
rect 27636 12236 27646 12292
rect 28242 12236 28252 12292
rect 28308 12236 33068 12292
rect 33124 12236 33134 12292
rect 34262 12236 34300 12292
rect 34356 12236 34366 12292
rect 34486 12236 34524 12292
rect 34580 12236 34590 12292
rect 35074 12236 35084 12292
rect 35140 12236 35868 12292
rect 35924 12236 35934 12292
rect 36754 12236 36764 12292
rect 36820 12236 36988 12292
rect 37044 12236 37054 12292
rect 38658 12236 38668 12292
rect 38724 12236 40908 12292
rect 40964 12236 40974 12292
rect 6290 12124 6300 12180
rect 6356 12124 10388 12180
rect 10546 12124 10556 12180
rect 10612 12124 11004 12180
rect 11060 12124 11070 12180
rect 12002 12124 12012 12180
rect 12068 12124 12572 12180
rect 12628 12124 12638 12180
rect 13458 12124 13468 12180
rect 13524 12124 13580 12180
rect 13636 12124 13646 12180
rect 14466 12124 14476 12180
rect 14532 12124 14542 12180
rect 16818 12124 16828 12180
rect 16884 12124 16940 12180
rect 16996 12124 17006 12180
rect 18060 12124 18172 12180
rect 18228 12124 18238 12180
rect 18620 12124 18956 12180
rect 19012 12124 22652 12180
rect 22708 12124 22718 12180
rect 23650 12124 23660 12180
rect 23716 12124 25340 12180
rect 25396 12124 25406 12180
rect 29110 12124 29148 12180
rect 29204 12124 29214 12180
rect 29586 12124 29596 12180
rect 29652 12124 30380 12180
rect 30436 12124 30446 12180
rect 30930 12124 30940 12180
rect 30996 12124 31164 12180
rect 31220 12124 31230 12180
rect 33842 12124 33852 12180
rect 33908 12124 34860 12180
rect 34916 12124 35308 12180
rect 35364 12124 35374 12180
rect 37650 12124 37660 12180
rect 37716 12124 40460 12180
rect 40516 12124 40526 12180
rect 9762 12012 9772 12068
rect 9828 12012 15820 12068
rect 15876 12012 15886 12068
rect 18060 11956 18116 12124
rect 18274 12012 18284 12068
rect 18340 12012 19404 12068
rect 19460 12012 19470 12068
rect 30482 12012 30492 12068
rect 30548 12012 30660 12068
rect 30790 12012 30828 12068
rect 30884 12012 30894 12068
rect 31042 12012 31052 12068
rect 31108 12012 31146 12068
rect 31490 12012 31500 12068
rect 31556 12012 33964 12068
rect 34020 12012 34030 12068
rect 34290 12012 34300 12068
rect 34356 12012 35756 12068
rect 35812 12012 35822 12068
rect 37426 12012 37436 12068
rect 37492 12012 38556 12068
rect 38612 12012 38622 12068
rect 38770 12012 38780 12068
rect 38836 12012 41916 12068
rect 41972 12012 41982 12068
rect 2818 11900 2828 11956
rect 2884 11900 4284 11956
rect 4340 11900 4900 11956
rect 5842 11900 5852 11956
rect 5908 11900 13692 11956
rect 13748 11900 13758 11956
rect 15586 11900 15596 11956
rect 15652 11900 19628 11956
rect 19684 11900 19694 11956
rect 20972 11900 27132 11956
rect 27188 11900 27916 11956
rect 27972 11900 27982 11956
rect 28242 11900 28252 11956
rect 28308 11900 28476 11956
rect 28532 11900 28542 11956
rect 4844 11844 4900 11900
rect 15820 11844 15876 11900
rect 20972 11844 21028 11900
rect 4844 11788 7196 11844
rect 7252 11788 8204 11844
rect 8260 11788 8652 11844
rect 8708 11788 9660 11844
rect 9716 11788 9726 11844
rect 10556 11788 11116 11844
rect 11172 11788 11182 11844
rect 11442 11788 11452 11844
rect 11508 11788 12348 11844
rect 12404 11788 12414 11844
rect 15250 11788 15260 11844
rect 15316 11788 15652 11844
rect 15810 11788 15820 11844
rect 15876 11788 15886 11844
rect 16034 11788 16044 11844
rect 16100 11788 17724 11844
rect 17780 11788 17790 11844
rect 20178 11788 20188 11844
rect 20244 11788 20972 11844
rect 21028 11788 21038 11844
rect 23538 11788 23548 11844
rect 23604 11788 24332 11844
rect 24388 11788 24398 11844
rect 30604 11788 30660 12012
rect 31154 11900 31164 11956
rect 31220 11900 31258 11956
rect 34178 11900 34188 11956
rect 34244 11900 38108 11956
rect 38164 11900 38174 11956
rect 32274 11788 32284 11844
rect 32340 11788 34412 11844
rect 34468 11788 34478 11844
rect 37426 11788 37436 11844
rect 37492 11788 38668 11844
rect 38724 11788 38734 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 10556 11732 10612 11788
rect 15596 11732 15652 11788
rect 30594 11732 30604 11788
rect 30660 11732 30670 11788
rect 31154 11732 31164 11788
rect 31220 11732 31258 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 10546 11676 10556 11732
rect 10612 11676 10622 11732
rect 11778 11676 11788 11732
rect 11844 11676 12460 11732
rect 12516 11676 12526 11732
rect 12758 11676 12796 11732
rect 12852 11676 12862 11732
rect 13794 11676 13804 11732
rect 13860 11676 14700 11732
rect 14756 11676 15148 11732
rect 15586 11676 15596 11732
rect 15652 11676 15662 11732
rect 16706 11676 16716 11732
rect 16772 11676 21756 11732
rect 21812 11676 23884 11732
rect 23940 11676 26908 11732
rect 26964 11676 27468 11732
rect 27524 11676 27534 11732
rect 29698 11676 29708 11732
rect 29764 11676 30044 11732
rect 30100 11676 30110 11732
rect 32946 11676 32956 11732
rect 33012 11676 34524 11732
rect 34580 11676 34590 11732
rect 35532 11676 37324 11732
rect 37380 11676 37390 11732
rect 37538 11676 37548 11732
rect 37604 11676 40068 11732
rect 11666 11564 11676 11620
rect 11732 11564 11742 11620
rect 11676 11508 11732 11564
rect 15092 11508 15148 11676
rect 35532 11620 35588 11676
rect 40012 11620 40068 11676
rect 15922 11564 15932 11620
rect 15988 11564 16604 11620
rect 16660 11564 16670 11620
rect 17042 11564 17052 11620
rect 17108 11564 22092 11620
rect 22148 11564 22876 11620
rect 22932 11564 22942 11620
rect 26674 11564 26684 11620
rect 26740 11564 26908 11620
rect 26964 11564 33740 11620
rect 33796 11564 33806 11620
rect 33964 11564 35588 11620
rect 35746 11564 35756 11620
rect 35812 11564 36092 11620
rect 36148 11564 38892 11620
rect 38948 11564 38958 11620
rect 40002 11564 40012 11620
rect 40068 11564 40460 11620
rect 40516 11564 40526 11620
rect 33964 11508 34020 11564
rect 10098 11452 10108 11508
rect 10164 11452 11732 11508
rect 12898 11452 12908 11508
rect 12964 11452 12974 11508
rect 13878 11452 13916 11508
rect 13972 11452 13982 11508
rect 15092 11452 16604 11508
rect 16660 11452 16670 11508
rect 19506 11452 19516 11508
rect 19572 11452 23212 11508
rect 23268 11452 23278 11508
rect 25442 11452 25452 11508
rect 25508 11452 25900 11508
rect 25956 11452 28700 11508
rect 28756 11452 28766 11508
rect 28914 11452 28924 11508
rect 28980 11452 32732 11508
rect 32788 11452 34020 11508
rect 34402 11452 34412 11508
rect 34468 11452 36764 11508
rect 36820 11452 36830 11508
rect 37090 11452 37100 11508
rect 37156 11452 37324 11508
rect 37380 11452 37772 11508
rect 37828 11452 37838 11508
rect 38658 11452 38668 11508
rect 38724 11452 40236 11508
rect 40292 11452 40302 11508
rect 12908 11396 12964 11452
rect 5292 11340 8092 11396
rect 8148 11340 8428 11396
rect 8484 11340 12124 11396
rect 12180 11340 13244 11396
rect 13300 11340 13310 11396
rect 14466 11340 14476 11396
rect 14532 11340 15932 11396
rect 15988 11340 15998 11396
rect 18834 11340 18844 11396
rect 18900 11340 19964 11396
rect 20020 11340 20030 11396
rect 25778 11340 25788 11396
rect 25844 11340 31164 11396
rect 31220 11340 31230 11396
rect 32806 11340 32844 11396
rect 32900 11340 32910 11396
rect 33170 11340 33180 11396
rect 33236 11340 39452 11396
rect 39508 11340 39518 11396
rect 39750 11340 39788 11396
rect 39844 11340 39854 11396
rect 5292 11172 5348 11340
rect 6066 11228 6076 11284
rect 6132 11228 8652 11284
rect 8708 11228 8718 11284
rect 10882 11228 10892 11284
rect 10948 11228 11676 11284
rect 11732 11228 11742 11284
rect 13346 11228 13356 11284
rect 13412 11228 14700 11284
rect 14756 11228 14766 11284
rect 16930 11228 16940 11284
rect 16996 11228 17276 11284
rect 17332 11228 17342 11284
rect 18386 11228 18396 11284
rect 18452 11228 27244 11284
rect 27300 11228 27310 11284
rect 27906 11228 27916 11284
rect 27972 11228 33516 11284
rect 33572 11228 33582 11284
rect 34178 11228 34188 11284
rect 34244 11228 34300 11284
rect 34356 11228 34636 11284
rect 34692 11228 34702 11284
rect 36754 11228 36764 11284
rect 36820 11228 37212 11284
rect 37268 11228 37660 11284
rect 37716 11228 37726 11284
rect 37874 11228 37884 11284
rect 37940 11228 38444 11284
rect 38500 11228 38510 11284
rect 39106 11228 39116 11284
rect 39172 11228 40460 11284
rect 40516 11228 40526 11284
rect 41234 11228 41244 11284
rect 41300 11228 42140 11284
rect 42196 11228 42206 11284
rect 3602 11116 3612 11172
rect 3668 11116 4060 11172
rect 4116 11116 4126 11172
rect 4498 11116 4508 11172
rect 4564 11116 5292 11172
rect 5348 11116 5358 11172
rect 6178 11116 6188 11172
rect 6244 11116 6748 11172
rect 6804 11116 9884 11172
rect 9940 11116 9950 11172
rect 10322 11116 10332 11172
rect 10388 11116 11004 11172
rect 11060 11116 11900 11172
rect 11956 11116 11966 11172
rect 13906 11116 13916 11172
rect 13972 11116 14476 11172
rect 14532 11116 14542 11172
rect 16818 11116 16828 11172
rect 16884 11116 20524 11172
rect 20580 11116 20590 11172
rect 22194 11116 22204 11172
rect 22260 11116 29652 11172
rect 29810 11116 29820 11172
rect 29876 11116 30828 11172
rect 30884 11116 36652 11172
rect 36708 11116 36718 11172
rect 37398 11116 37436 11172
rect 37492 11116 37502 11172
rect 37650 11116 37660 11172
rect 37716 11116 38668 11172
rect 38882 11116 38892 11172
rect 38948 11116 40572 11172
rect 40628 11116 41692 11172
rect 41748 11116 41758 11172
rect 29596 11060 29652 11116
rect 38612 11060 38668 11116
rect 4946 11004 4956 11060
rect 5012 11004 6972 11060
rect 7028 11004 7644 11060
rect 7700 11004 7710 11060
rect 7858 11004 7868 11060
rect 7924 11004 8876 11060
rect 8932 11004 8942 11060
rect 15362 11004 15372 11060
rect 15428 11004 18004 11060
rect 22866 11004 22876 11060
rect 22932 11004 27580 11060
rect 27636 11004 28700 11060
rect 28756 11004 28766 11060
rect 29596 11004 30044 11060
rect 30100 11004 30110 11060
rect 32274 11004 32284 11060
rect 32340 11004 36092 11060
rect 36148 11004 38444 11060
rect 38500 11004 38510 11060
rect 38612 11004 38892 11060
rect 38948 11004 38958 11060
rect 39778 11004 39788 11060
rect 39844 11004 40236 11060
rect 40292 11004 40302 11060
rect 7644 10948 7700 11004
rect 17948 10948 18004 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 7644 10892 8988 10948
rect 9044 10892 9054 10948
rect 13906 10892 13916 10948
rect 13972 10892 17724 10948
rect 17780 10892 17790 10948
rect 17938 10892 17948 10948
rect 18004 10892 19012 10948
rect 19478 10892 19516 10948
rect 19572 10892 19582 10948
rect 28354 10892 28364 10948
rect 28420 10892 29708 10948
rect 29764 10892 29774 10948
rect 31378 10892 31388 10948
rect 31444 10892 31836 10948
rect 31892 10892 34076 10948
rect 34132 10892 34636 10948
rect 34692 10892 34860 10948
rect 34916 10892 35532 10948
rect 35588 10892 35598 10948
rect 35970 10892 35980 10948
rect 36036 10892 36316 10948
rect 36372 10892 36382 10948
rect 37660 10892 40348 10948
rect 40404 10892 40414 10948
rect 18956 10836 19012 10892
rect 2706 10780 2716 10836
rect 2772 10780 5180 10836
rect 5236 10780 5246 10836
rect 12450 10780 12460 10836
rect 12516 10780 13020 10836
rect 13076 10780 13086 10836
rect 18274 10780 18284 10836
rect 18340 10780 18732 10836
rect 18788 10780 18798 10836
rect 18956 10780 20076 10836
rect 20132 10780 22204 10836
rect 22260 10780 22270 10836
rect 24630 10780 24668 10836
rect 24724 10780 24734 10836
rect 26114 10780 26124 10836
rect 26180 10780 27916 10836
rect 27972 10780 29148 10836
rect 29204 10780 29214 10836
rect 32610 10780 32620 10836
rect 32676 10780 34300 10836
rect 34356 10780 34366 10836
rect 34626 10780 34636 10836
rect 34692 10780 34972 10836
rect 35028 10780 35038 10836
rect 35970 10780 35980 10836
rect 36036 10780 36428 10836
rect 36484 10780 36494 10836
rect 6290 10668 6300 10724
rect 6356 10668 9884 10724
rect 9940 10668 12908 10724
rect 12964 10668 12974 10724
rect 16482 10668 16492 10724
rect 16548 10668 17612 10724
rect 17668 10668 17678 10724
rect 18162 10668 18172 10724
rect 18228 10668 19068 10724
rect 19124 10668 19516 10724
rect 19572 10668 20188 10724
rect 20244 10668 20254 10724
rect 23426 10668 23436 10724
rect 23492 10668 25900 10724
rect 25956 10668 25966 10724
rect 26562 10668 26572 10724
rect 26628 10668 28364 10724
rect 28420 10668 31388 10724
rect 31444 10668 31454 10724
rect 33730 10668 33740 10724
rect 33796 10668 36540 10724
rect 36596 10668 36606 10724
rect 37660 10612 37716 10892
rect 38434 10780 38444 10836
rect 38500 10780 38668 10836
rect 39554 10780 39564 10836
rect 39620 10780 41692 10836
rect 41748 10780 41758 10836
rect 38612 10724 38668 10780
rect 38612 10668 39732 10724
rect 6850 10556 6860 10612
rect 6916 10556 8316 10612
rect 8372 10556 8382 10612
rect 16594 10556 16604 10612
rect 16660 10556 19964 10612
rect 20020 10556 20030 10612
rect 26852 10556 28028 10612
rect 28084 10556 31500 10612
rect 31556 10556 33628 10612
rect 33684 10556 33694 10612
rect 34514 10556 34524 10612
rect 34580 10556 34972 10612
rect 35028 10556 35038 10612
rect 35298 10556 35308 10612
rect 35364 10556 35980 10612
rect 36036 10556 36046 10612
rect 37426 10556 37436 10612
rect 37492 10556 37502 10612
rect 37650 10556 37660 10612
rect 37716 10556 37726 10612
rect 26852 10500 26908 10556
rect 37436 10500 37492 10556
rect 39676 10500 39732 10668
rect 4050 10444 4060 10500
rect 4116 10444 5740 10500
rect 5796 10444 9996 10500
rect 10052 10444 10062 10500
rect 17462 10444 17500 10500
rect 17556 10444 17566 10500
rect 25666 10444 25676 10500
rect 25732 10444 25900 10500
rect 25956 10444 26908 10500
rect 32498 10444 32508 10500
rect 32564 10444 37100 10500
rect 37156 10444 37166 10500
rect 37436 10444 38220 10500
rect 38276 10444 38286 10500
rect 39676 10444 40460 10500
rect 40516 10444 40526 10500
rect 4274 10332 4284 10388
rect 4340 10332 9884 10388
rect 9940 10332 9950 10388
rect 16594 10332 16604 10388
rect 16660 10332 18172 10388
rect 18228 10332 18732 10388
rect 18788 10332 18798 10388
rect 23650 10332 23660 10388
rect 23716 10332 24444 10388
rect 24500 10332 25452 10388
rect 25508 10332 26012 10388
rect 26068 10332 26078 10388
rect 28690 10332 28700 10388
rect 28756 10332 32732 10388
rect 32788 10332 32798 10388
rect 32956 10332 33292 10388
rect 33348 10332 35308 10388
rect 35364 10332 35374 10388
rect 36082 10332 36092 10388
rect 36148 10332 36428 10388
rect 36484 10332 36494 10388
rect 36642 10332 36652 10388
rect 36708 10332 36764 10388
rect 36820 10332 36830 10388
rect 39330 10332 39340 10388
rect 39396 10332 41692 10388
rect 41748 10332 41758 10388
rect 32956 10276 33012 10332
rect 17602 10220 17612 10276
rect 17668 10220 17724 10276
rect 17780 10220 17790 10276
rect 22754 10220 22764 10276
rect 22820 10220 26796 10276
rect 26852 10220 26862 10276
rect 31378 10220 31388 10276
rect 31444 10220 33012 10276
rect 36530 10220 36540 10276
rect 36596 10220 37100 10276
rect 37156 10220 37166 10276
rect 37426 10220 37436 10276
rect 37492 10220 43260 10276
rect 43316 10220 43326 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 16594 10108 16604 10164
rect 16660 10108 21980 10164
rect 22036 10108 22046 10164
rect 24994 10108 25004 10164
rect 25060 10108 25564 10164
rect 25620 10108 25630 10164
rect 26338 10108 26348 10164
rect 26404 10108 27804 10164
rect 27860 10108 27870 10164
rect 29810 10108 29820 10164
rect 29876 10108 32844 10164
rect 32900 10108 32910 10164
rect 34262 10108 34300 10164
rect 34356 10108 34366 10164
rect 34598 10108 34636 10164
rect 34692 10108 34702 10164
rect 35970 10108 35980 10164
rect 36036 10108 38220 10164
rect 38276 10108 38286 10164
rect 39778 10108 39788 10164
rect 39844 10108 40908 10164
rect 40964 10108 41188 10164
rect 41132 10052 41188 10108
rect 3266 9996 3276 10052
rect 3332 9996 3612 10052
rect 3668 9996 4508 10052
rect 4564 9996 5628 10052
rect 5684 9996 5694 10052
rect 6738 9996 6748 10052
rect 6804 9996 7420 10052
rect 7476 9996 7486 10052
rect 17490 9996 17500 10052
rect 17556 9996 17566 10052
rect 17714 9996 17724 10052
rect 17780 9996 18396 10052
rect 18452 9996 18462 10052
rect 19170 9996 19180 10052
rect 19236 9996 20860 10052
rect 20916 9996 21644 10052
rect 21700 9996 21710 10052
rect 22278 9996 22316 10052
rect 22372 9996 22382 10052
rect 25666 9996 25676 10052
rect 25732 9996 26684 10052
rect 26740 9996 26750 10052
rect 28914 9996 28924 10052
rect 28980 9996 29596 10052
rect 29652 9996 29662 10052
rect 30258 9996 30268 10052
rect 30324 9996 33964 10052
rect 34020 9996 35868 10052
rect 35924 9996 35934 10052
rect 37762 9996 37772 10052
rect 37828 9996 39620 10052
rect 40338 9996 40348 10052
rect 40404 9996 40796 10052
rect 40852 9996 40862 10052
rect 41132 9996 41468 10052
rect 41524 9996 41534 10052
rect 17500 9940 17556 9996
rect 35868 9940 35924 9996
rect 39564 9940 39620 9996
rect 5058 9884 5068 9940
rect 5124 9884 5964 9940
rect 6020 9884 8988 9940
rect 9044 9884 9436 9940
rect 9492 9884 9772 9940
rect 9828 9884 11900 9940
rect 11956 9884 13804 9940
rect 13860 9884 13870 9940
rect 17500 9884 19404 9940
rect 19460 9884 19470 9940
rect 20738 9884 20748 9940
rect 20804 9884 22540 9940
rect 22596 9884 22606 9940
rect 27682 9884 27692 9940
rect 27748 9884 29484 9940
rect 29540 9884 30044 9940
rect 30100 9884 30110 9940
rect 30594 9884 30604 9940
rect 30660 9884 31164 9940
rect 31220 9884 31230 9940
rect 35298 9884 35308 9940
rect 35364 9884 35644 9940
rect 35700 9884 35710 9940
rect 35868 9884 37884 9940
rect 37940 9884 37950 9940
rect 39554 9884 39564 9940
rect 39620 9884 41076 9940
rect 3826 9772 3836 9828
rect 3892 9772 10108 9828
rect 10164 9772 10174 9828
rect 11554 9772 11564 9828
rect 11620 9772 13132 9828
rect 13188 9772 13198 9828
rect 17490 9772 17500 9828
rect 17556 9772 19068 9828
rect 19124 9772 19134 9828
rect 22082 9772 22092 9828
rect 22148 9772 22316 9828
rect 22372 9772 22382 9828
rect 23202 9772 23212 9828
rect 23268 9772 23772 9828
rect 23828 9772 26908 9828
rect 27346 9772 27356 9828
rect 27412 9772 28140 9828
rect 28196 9772 29372 9828
rect 29428 9772 29438 9828
rect 29586 9772 29596 9828
rect 29652 9772 31612 9828
rect 31668 9772 31678 9828
rect 36082 9772 36092 9828
rect 36148 9772 36204 9828
rect 36260 9772 36270 9828
rect 37538 9772 37548 9828
rect 37604 9772 38556 9828
rect 4834 9660 4844 9716
rect 4900 9660 6076 9716
rect 6132 9660 9212 9716
rect 9268 9660 9278 9716
rect 10882 9660 10892 9716
rect 10948 9660 12796 9716
rect 12852 9660 13916 9716
rect 13972 9660 13982 9716
rect 14130 9660 14140 9716
rect 14196 9660 17724 9716
rect 17780 9660 17790 9716
rect 18834 9660 18844 9716
rect 18900 9660 19180 9716
rect 19236 9660 19246 9716
rect 23986 9660 23996 9716
rect 24052 9660 25564 9716
rect 25620 9660 25630 9716
rect 26852 9604 26908 9772
rect 38612 9716 38668 9828
rect 38770 9772 38780 9828
rect 38836 9772 40348 9828
rect 40404 9772 40414 9828
rect 40674 9772 40684 9828
rect 40740 9772 40796 9828
rect 40852 9772 40862 9828
rect 27458 9660 27468 9716
rect 27524 9660 28812 9716
rect 28868 9660 28878 9716
rect 30818 9660 30828 9716
rect 30884 9660 37436 9716
rect 37492 9660 37502 9716
rect 38612 9660 40572 9716
rect 40628 9660 40638 9716
rect 41020 9604 41076 9884
rect 41906 9772 41916 9828
rect 41972 9772 41982 9828
rect 41570 9660 41580 9716
rect 41636 9660 41692 9716
rect 41748 9660 41758 9716
rect 3332 9548 3836 9604
rect 3892 9548 3902 9604
rect 4162 9548 4172 9604
rect 4228 9548 7644 9604
rect 7700 9548 7710 9604
rect 13794 9548 13804 9604
rect 13860 9548 16828 9604
rect 16884 9548 18396 9604
rect 18452 9548 18462 9604
rect 18610 9548 18620 9604
rect 18676 9548 26684 9604
rect 26740 9548 26750 9604
rect 26852 9548 28588 9604
rect 28644 9548 28654 9604
rect 30146 9548 30156 9604
rect 30212 9548 31052 9604
rect 31108 9548 31118 9604
rect 31266 9548 31276 9604
rect 31332 9548 31948 9604
rect 32004 9548 36260 9604
rect 38770 9548 38780 9604
rect 38836 9548 39788 9604
rect 39844 9548 39854 9604
rect 40898 9548 40908 9604
rect 40964 9548 41356 9604
rect 41412 9548 41422 9604
rect 3332 9492 3388 9548
rect 1810 9436 1820 9492
rect 1876 9436 3388 9492
rect 3602 9436 3612 9492
rect 3668 9436 7196 9492
rect 7252 9436 7262 9492
rect 18274 9436 18284 9492
rect 18340 9436 19516 9492
rect 19572 9436 19582 9492
rect 22978 9436 22988 9492
rect 23044 9436 26460 9492
rect 26516 9436 26526 9492
rect 3612 9380 3668 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 26684 9380 26740 9548
rect 28588 9492 28644 9548
rect 28588 9436 32060 9492
rect 32116 9436 32126 9492
rect 33506 9436 33516 9492
rect 33572 9436 35980 9492
rect 36036 9436 36046 9492
rect 36204 9380 36260 9548
rect 41916 9492 41972 9772
rect 36978 9436 36988 9492
rect 37044 9436 37324 9492
rect 37380 9436 37390 9492
rect 37650 9436 37660 9492
rect 37716 9436 39004 9492
rect 39060 9436 39070 9492
rect 39218 9436 39228 9492
rect 39284 9436 39564 9492
rect 39620 9436 39676 9492
rect 39732 9436 39742 9492
rect 39890 9436 39900 9492
rect 39956 9436 41972 9492
rect 2594 9324 2604 9380
rect 2660 9324 3668 9380
rect 4386 9324 4396 9380
rect 4452 9324 5740 9380
rect 5796 9324 9156 9380
rect 17574 9324 17612 9380
rect 17668 9324 17678 9380
rect 22418 9324 22428 9380
rect 22484 9324 23996 9380
rect 24052 9324 24062 9380
rect 24546 9324 24556 9380
rect 24612 9324 25676 9380
rect 25732 9324 25742 9380
rect 26674 9324 26684 9380
rect 26740 9324 26750 9380
rect 27122 9324 27132 9380
rect 27188 9324 33740 9380
rect 33796 9324 33806 9380
rect 35522 9324 35532 9380
rect 35588 9324 35868 9380
rect 35924 9324 35934 9380
rect 36204 9324 39788 9380
rect 39844 9324 39854 9380
rect 9100 9268 9156 9324
rect 5254 9212 5292 9268
rect 5348 9212 5358 9268
rect 7970 9212 7980 9268
rect 8036 9212 8764 9268
rect 8820 9212 8830 9268
rect 9090 9212 9100 9268
rect 9156 9212 9884 9268
rect 9940 9212 10780 9268
rect 10836 9212 10846 9268
rect 17042 9212 17052 9268
rect 17108 9212 17724 9268
rect 17780 9212 17790 9268
rect 23538 9212 23548 9268
rect 23604 9212 27244 9268
rect 27300 9212 27310 9268
rect 28364 9212 28476 9268
rect 28532 9212 28542 9268
rect 29026 9212 29036 9268
rect 29092 9212 29260 9268
rect 29316 9212 29596 9268
rect 29652 9212 29662 9268
rect 32162 9212 32172 9268
rect 32228 9212 33852 9268
rect 33908 9212 33918 9268
rect 34076 9212 39228 9268
rect 39284 9212 39294 9268
rect 39442 9212 39452 9268
rect 39508 9212 39676 9268
rect 39732 9212 39742 9268
rect 41794 9212 41804 9268
rect 41860 9212 41916 9268
rect 41972 9212 41982 9268
rect 1922 9100 1932 9156
rect 1988 9100 3724 9156
rect 3780 9100 4844 9156
rect 4900 9100 4910 9156
rect 5394 9100 5404 9156
rect 5460 9100 6076 9156
rect 6132 9100 6142 9156
rect 7074 9100 7084 9156
rect 7140 9100 8876 9156
rect 8932 9100 8942 9156
rect 10098 9100 10108 9156
rect 10164 9100 12012 9156
rect 12068 9100 12572 9156
rect 12628 9100 12638 9156
rect 17042 9100 17052 9156
rect 17108 9100 18508 9156
rect 18564 9100 18956 9156
rect 19012 9100 19022 9156
rect 22306 9100 22316 9156
rect 22372 9100 24668 9156
rect 24724 9100 24734 9156
rect 26086 9100 26124 9156
rect 26180 9100 26190 9156
rect 26450 9100 26460 9156
rect 26516 9100 27804 9156
rect 27860 9100 27870 9156
rect 26124 9044 26180 9100
rect 28364 9044 28420 9212
rect 34076 9156 34132 9212
rect 28578 9100 28588 9156
rect 28644 9100 34132 9156
rect 34524 9100 36428 9156
rect 36484 9100 36494 9156
rect 36642 9100 36652 9156
rect 36708 9100 40572 9156
rect 40628 9100 41692 9156
rect 41748 9100 41758 9156
rect 3332 8988 5180 9044
rect 5236 8988 5246 9044
rect 6290 8988 6300 9044
rect 6356 8988 7308 9044
rect 7364 8988 7756 9044
rect 7812 8988 10220 9044
rect 10276 8988 10286 9044
rect 19506 8988 19516 9044
rect 19572 8988 22540 9044
rect 22596 8988 22988 9044
rect 23044 8988 23054 9044
rect 23538 8988 23548 9044
rect 23604 8988 24108 9044
rect 24164 8988 24174 9044
rect 24770 8988 24780 9044
rect 24836 8988 26180 9044
rect 27906 8988 27916 9044
rect 27972 8988 31164 9044
rect 31220 8988 31230 9044
rect 31378 8988 31388 9044
rect 31444 8988 32284 9044
rect 32340 8988 32350 9044
rect 3332 8932 3388 8988
rect 34524 8932 34580 9100
rect 34672 8988 34748 9044
rect 34804 8988 37996 9044
rect 38052 8988 38062 9044
rect 38210 8988 38220 9044
rect 38276 8988 39676 9044
rect 39732 8988 39742 9044
rect 40450 8988 40460 9044
rect 40516 8988 40796 9044
rect 40852 8988 40862 9044
rect 3042 8876 3052 8932
rect 3108 8876 3388 8932
rect 4050 8876 4060 8932
rect 4116 8876 4284 8932
rect 4340 8876 4350 8932
rect 6850 8876 6860 8932
rect 6916 8876 8092 8932
rect 8148 8876 8158 8932
rect 8978 8876 8988 8932
rect 9044 8876 10556 8932
rect 10612 8876 10622 8932
rect 17266 8876 17276 8932
rect 17332 8876 18172 8932
rect 18228 8876 18238 8932
rect 18834 8876 18844 8932
rect 18900 8876 19180 8932
rect 19236 8876 21644 8932
rect 21700 8876 21710 8932
rect 23090 8876 23100 8932
rect 23156 8876 23660 8932
rect 23716 8876 23726 8932
rect 25666 8876 25676 8932
rect 25732 8876 28252 8932
rect 28308 8876 28318 8932
rect 29586 8876 29596 8932
rect 29652 8876 34580 8932
rect 34850 8876 34860 8932
rect 34916 8876 35532 8932
rect 35588 8876 36876 8932
rect 36932 8876 36942 8932
rect 39778 8876 39788 8932
rect 39844 8876 42140 8932
rect 42196 8876 42206 8932
rect 21644 8820 21700 8876
rect 3490 8764 3500 8820
rect 3556 8764 7252 8820
rect 7410 8764 7420 8820
rect 7476 8764 8652 8820
rect 8708 8764 8718 8820
rect 8866 8764 8876 8820
rect 8932 8764 9212 8820
rect 9268 8764 11564 8820
rect 11620 8764 11630 8820
rect 21644 8764 24220 8820
rect 24276 8764 24286 8820
rect 24658 8764 24668 8820
rect 24724 8764 26236 8820
rect 26292 8764 26302 8820
rect 34962 8764 34972 8820
rect 35028 8764 35420 8820
rect 35476 8764 37156 8820
rect 37286 8764 37324 8820
rect 37380 8764 37390 8820
rect 39330 8764 39340 8820
rect 39396 8764 41356 8820
rect 41412 8764 41422 8820
rect 7196 8708 7252 8764
rect 37100 8708 37156 8764
rect 7196 8652 9772 8708
rect 9828 8652 17388 8708
rect 17444 8652 17454 8708
rect 17938 8652 17948 8708
rect 18004 8652 19180 8708
rect 19236 8652 19246 8708
rect 24322 8652 24332 8708
rect 24388 8652 25788 8708
rect 25844 8652 25854 8708
rect 37100 8652 37660 8708
rect 37716 8652 37726 8708
rect 38098 8652 38108 8708
rect 38164 8652 38444 8708
rect 38500 8652 38510 8708
rect 40338 8652 40348 8708
rect 40404 8652 41244 8708
rect 41300 8652 41310 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 38108 8596 38164 8652
rect 5058 8540 5068 8596
rect 5124 8540 5964 8596
rect 6020 8540 6030 8596
rect 7746 8540 7756 8596
rect 7812 8540 11676 8596
rect 11732 8540 11742 8596
rect 24630 8540 24668 8596
rect 24724 8540 24734 8596
rect 26786 8540 26796 8596
rect 26852 8540 28364 8596
rect 28420 8540 28430 8596
rect 29026 8540 29036 8596
rect 29092 8540 29484 8596
rect 29540 8540 29550 8596
rect 31714 8540 31724 8596
rect 31780 8540 33628 8596
rect 33684 8540 33694 8596
rect 36418 8540 36428 8596
rect 36484 8540 38164 8596
rect 39330 8540 39340 8596
rect 39396 8540 41020 8596
rect 41076 8540 41086 8596
rect 4946 8428 4956 8484
rect 5012 8428 5292 8484
rect 5348 8428 8652 8484
rect 8708 8428 8718 8484
rect 10294 8428 10332 8484
rect 10388 8428 10398 8484
rect 15250 8428 15260 8484
rect 15316 8428 15596 8484
rect 15652 8428 15662 8484
rect 18386 8428 18396 8484
rect 18452 8428 20524 8484
rect 20580 8428 21196 8484
rect 21252 8428 23548 8484
rect 23604 8428 23614 8484
rect 32050 8428 32060 8484
rect 32116 8428 38388 8484
rect 38658 8428 38668 8484
rect 38724 8428 39004 8484
rect 39060 8428 42476 8484
rect 42532 8428 42542 8484
rect 2146 8316 2156 8372
rect 2212 8316 3164 8372
rect 3220 8316 3230 8372
rect 4722 8316 4732 8372
rect 4788 8316 5068 8372
rect 5124 8316 5134 8372
rect 5394 8316 5404 8372
rect 5460 8316 5628 8372
rect 5684 8316 8204 8372
rect 8260 8316 9436 8372
rect 9492 8316 10892 8372
rect 10948 8316 10958 8372
rect 11442 8316 11452 8372
rect 11508 8316 12124 8372
rect 12180 8316 12190 8372
rect 15138 8316 15148 8372
rect 15204 8316 15708 8372
rect 15764 8316 15774 8372
rect 18050 8316 18060 8372
rect 18116 8316 20860 8372
rect 20916 8316 22428 8372
rect 22484 8316 22876 8372
rect 22932 8316 25228 8372
rect 25284 8316 25294 8372
rect 29362 8316 29372 8372
rect 29428 8316 29596 8372
rect 29652 8316 29662 8372
rect 30482 8316 30492 8372
rect 30548 8316 31388 8372
rect 31444 8316 31454 8372
rect 33394 8316 33404 8372
rect 33460 8316 36428 8372
rect 36484 8316 36494 8372
rect 38332 8260 38388 8428
rect 39554 8316 39564 8372
rect 39620 8316 40348 8372
rect 40404 8316 40684 8372
rect 40740 8316 40750 8372
rect 1922 8204 1932 8260
rect 1988 8204 3052 8260
rect 3108 8204 4172 8260
rect 4228 8204 4844 8260
rect 4900 8204 9660 8260
rect 9716 8204 9726 8260
rect 10658 8204 10668 8260
rect 10724 8204 11340 8260
rect 11396 8204 11406 8260
rect 12226 8204 12236 8260
rect 12292 8204 12460 8260
rect 12516 8204 12526 8260
rect 14018 8204 14028 8260
rect 14084 8204 14812 8260
rect 14868 8204 14878 8260
rect 15026 8204 15036 8260
rect 15092 8204 19964 8260
rect 20020 8204 20030 8260
rect 26114 8204 26124 8260
rect 26180 8204 35644 8260
rect 35700 8204 35710 8260
rect 36278 8204 36316 8260
rect 36372 8204 36382 8260
rect 38070 8204 38108 8260
rect 38164 8204 38174 8260
rect 38322 8204 38332 8260
rect 38388 8204 38398 8260
rect 10668 8148 10724 8204
rect 5618 8092 5628 8148
rect 5684 8092 6692 8148
rect 7186 8092 7196 8148
rect 7252 8092 7588 8148
rect 7858 8092 7868 8148
rect 7924 8092 10724 8148
rect 5628 8036 5684 8092
rect 6636 8036 6692 8092
rect 7532 8036 7588 8092
rect 12236 8036 12292 8204
rect 21298 8092 21308 8148
rect 21364 8092 29372 8148
rect 29428 8092 29438 8148
rect 35756 8092 37772 8148
rect 37828 8092 37838 8148
rect 39666 8092 39676 8148
rect 39732 8092 41020 8148
rect 41076 8092 41468 8148
rect 41524 8092 41534 8148
rect 41682 8092 41692 8148
rect 41748 8092 41786 8148
rect 35756 8036 35812 8092
rect 2146 7980 2156 8036
rect 2212 7980 2828 8036
rect 2884 7980 5012 8036
rect 5170 7980 5180 8036
rect 5236 7980 5684 8036
rect 5814 7980 5852 8036
rect 5908 7980 5918 8036
rect 6626 7980 6636 8036
rect 6692 7980 7084 8036
rect 7140 7980 7150 8036
rect 7522 7980 7532 8036
rect 7588 7980 12292 8036
rect 19730 7980 19740 8036
rect 19796 7980 21812 8036
rect 22082 7980 22092 8036
rect 22148 7980 23100 8036
rect 23156 7980 23166 8036
rect 26450 7980 26460 8036
rect 26516 7980 29708 8036
rect 29764 7980 29774 8036
rect 30566 7980 30604 8036
rect 30660 7980 33740 8036
rect 33796 7980 33806 8036
rect 35308 7980 35756 8036
rect 35812 7980 35822 8036
rect 36306 7980 36316 8036
rect 36372 7980 37884 8036
rect 37940 7980 37950 8036
rect 38994 7980 39004 8036
rect 39060 7980 39788 8036
rect 39844 7980 39854 8036
rect 40226 7980 40236 8036
rect 40292 7980 41580 8036
rect 41636 7980 41646 8036
rect 4956 7924 5012 7980
rect 21756 7924 21812 7980
rect 35308 7924 35364 7980
rect 2258 7868 2268 7924
rect 2324 7868 4900 7924
rect 4956 7868 9100 7924
rect 9156 7868 16044 7924
rect 16100 7868 16110 7924
rect 21746 7868 21756 7924
rect 21812 7868 21822 7924
rect 21980 7868 28700 7924
rect 28756 7868 28766 7924
rect 30930 7868 30940 7924
rect 30996 7868 31612 7924
rect 31668 7868 33068 7924
rect 33124 7868 35364 7924
rect 35522 7868 35532 7924
rect 35588 7868 36092 7924
rect 36148 7868 36316 7924
rect 36372 7868 41804 7924
rect 41860 7868 41870 7924
rect 2594 7756 2604 7812
rect 2660 7756 4508 7812
rect 4564 7756 4574 7812
rect 4844 7700 4900 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 21980 7812 22036 7868
rect 5058 7756 5068 7812
rect 5124 7756 6748 7812
rect 6804 7756 6814 7812
rect 20514 7756 20524 7812
rect 20580 7756 21420 7812
rect 21476 7756 21980 7812
rect 22036 7756 22046 7812
rect 24780 7756 26908 7812
rect 26964 7756 27468 7812
rect 27524 7756 27534 7812
rect 30594 7756 30604 7812
rect 30660 7756 31276 7812
rect 31332 7756 31342 7812
rect 32498 7756 32508 7812
rect 32564 7756 33516 7812
rect 33572 7756 33628 7812
rect 33684 7756 33694 7812
rect 35410 7756 35420 7812
rect 35476 7756 35644 7812
rect 35700 7756 35710 7812
rect 36754 7756 36764 7812
rect 36820 7756 36988 7812
rect 37044 7756 37054 7812
rect 37314 7756 37324 7812
rect 37380 7756 38332 7812
rect 38388 7756 38398 7812
rect 38612 7756 38892 7812
rect 38948 7756 38958 7812
rect 40114 7756 40124 7812
rect 40180 7756 41916 7812
rect 41972 7756 41982 7812
rect 2706 7644 2716 7700
rect 2772 7644 3612 7700
rect 3668 7644 4620 7700
rect 4676 7644 4686 7700
rect 4844 7644 7420 7700
rect 7476 7644 9996 7700
rect 10052 7644 12236 7700
rect 12292 7644 12302 7700
rect 13458 7644 13468 7700
rect 13524 7644 14252 7700
rect 14308 7644 19852 7700
rect 19908 7644 19918 7700
rect 24780 7588 24836 7756
rect 38612 7700 38668 7756
rect 29362 7644 29372 7700
rect 29428 7644 29708 7700
rect 29764 7644 30492 7700
rect 30548 7644 30558 7700
rect 30706 7644 30716 7700
rect 30772 7644 38668 7700
rect 39106 7644 39116 7700
rect 39172 7644 39900 7700
rect 39956 7644 39966 7700
rect 41234 7644 41244 7700
rect 41300 7644 41692 7700
rect 41748 7644 41972 7700
rect 3714 7532 3724 7588
rect 3780 7532 6972 7588
rect 7028 7532 7038 7588
rect 8866 7532 8876 7588
rect 8932 7532 10108 7588
rect 10164 7532 10174 7588
rect 20626 7532 20636 7588
rect 20692 7532 24780 7588
rect 24836 7532 24846 7588
rect 27906 7532 27916 7588
rect 27972 7532 38668 7588
rect 38612 7476 38668 7532
rect 4386 7420 4396 7476
rect 4452 7420 10668 7476
rect 10724 7420 10734 7476
rect 23650 7420 23660 7476
rect 23716 7420 25788 7476
rect 25844 7420 25854 7476
rect 28130 7420 28140 7476
rect 28196 7420 28476 7476
rect 28532 7420 29428 7476
rect 29586 7420 29596 7476
rect 29652 7420 30492 7476
rect 30548 7420 30558 7476
rect 30818 7420 30828 7476
rect 30884 7420 33628 7476
rect 33684 7420 33694 7476
rect 34850 7420 34860 7476
rect 34916 7420 36764 7476
rect 36820 7420 36830 7476
rect 38612 7420 40684 7476
rect 40740 7420 40750 7476
rect 29372 7364 29428 7420
rect 41916 7364 41972 7644
rect 5142 7308 5180 7364
rect 5236 7308 5246 7364
rect 6850 7308 6860 7364
rect 6916 7308 8652 7364
rect 8708 7308 8718 7364
rect 9650 7308 9660 7364
rect 9716 7308 11788 7364
rect 11844 7308 12796 7364
rect 12852 7308 12862 7364
rect 18610 7308 18620 7364
rect 18676 7308 20636 7364
rect 20692 7308 20702 7364
rect 21298 7308 21308 7364
rect 21364 7308 24444 7364
rect 24500 7308 24892 7364
rect 24948 7308 24958 7364
rect 27682 7308 27692 7364
rect 27748 7308 28588 7364
rect 28644 7308 28654 7364
rect 28802 7308 28812 7364
rect 28868 7308 28878 7364
rect 29372 7308 30604 7364
rect 30660 7308 30670 7364
rect 34626 7308 34636 7364
rect 34692 7308 35308 7364
rect 35364 7308 36316 7364
rect 36372 7308 37268 7364
rect 41906 7308 41916 7364
rect 41972 7308 41982 7364
rect 28812 7252 28868 7308
rect 2482 7196 2492 7252
rect 2548 7196 5628 7252
rect 5684 7196 5694 7252
rect 5842 7196 5852 7252
rect 5908 7196 11116 7252
rect 11172 7196 11182 7252
rect 28736 7196 28812 7252
rect 28868 7196 30716 7252
rect 30772 7196 30782 7252
rect 32274 7196 32284 7252
rect 32340 7196 35084 7252
rect 35140 7196 36540 7252
rect 36596 7196 36606 7252
rect 37212 7140 37268 7308
rect 41346 7196 41356 7252
rect 41412 7196 41692 7252
rect 41748 7196 41758 7252
rect 4834 7084 4844 7140
rect 4900 7084 5292 7140
rect 5348 7084 5740 7140
rect 5796 7084 5806 7140
rect 6066 7084 6076 7140
rect 6132 7084 6524 7140
rect 6580 7084 6590 7140
rect 14018 7084 14028 7140
rect 14084 7084 20524 7140
rect 20580 7084 20590 7140
rect 23202 7084 23212 7140
rect 23268 7084 23996 7140
rect 24052 7084 27916 7140
rect 27972 7084 27982 7140
rect 28802 7084 28812 7140
rect 28868 7084 29260 7140
rect 29316 7084 29326 7140
rect 37202 7084 37212 7140
rect 37268 7084 37278 7140
rect 40674 7084 40684 7140
rect 40740 7084 42028 7140
rect 42084 7084 42094 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 23212 7028 23268 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 5282 6972 5292 7028
rect 5348 6972 6300 7028
rect 6356 6972 6366 7028
rect 16566 6972 16604 7028
rect 16660 6972 16670 7028
rect 18274 6972 18284 7028
rect 18340 6972 23268 7028
rect 24882 6972 24892 7028
rect 24948 6972 29932 7028
rect 29988 6972 29998 7028
rect 13458 6860 13468 6916
rect 13524 6860 17276 6916
rect 17332 6860 17342 6916
rect 26852 6860 29820 6916
rect 29876 6860 29886 6916
rect 39218 6860 39228 6916
rect 39284 6860 40572 6916
rect 40628 6860 41804 6916
rect 41860 6860 41870 6916
rect 26852 6804 26908 6860
rect 3602 6748 3612 6804
rect 3668 6748 6524 6804
rect 6580 6748 6590 6804
rect 9426 6748 9436 6804
rect 9492 6748 9660 6804
rect 9716 6748 9726 6804
rect 12786 6748 12796 6804
rect 12852 6748 13916 6804
rect 13972 6748 14252 6804
rect 14308 6748 16156 6804
rect 16212 6748 16222 6804
rect 19842 6748 19852 6804
rect 19908 6748 21420 6804
rect 21476 6748 21486 6804
rect 24658 6748 24668 6804
rect 24724 6748 24734 6804
rect 24994 6748 25004 6804
rect 25060 6748 26908 6804
rect 29922 6748 29932 6804
rect 29988 6748 40796 6804
rect 40852 6748 40862 6804
rect 3154 6636 3164 6692
rect 3220 6636 5292 6692
rect 5348 6636 5358 6692
rect 5964 6580 6020 6748
rect 24668 6692 24724 6748
rect 7746 6636 7756 6692
rect 7812 6636 9884 6692
rect 9940 6636 13020 6692
rect 13076 6636 13086 6692
rect 15362 6636 15372 6692
rect 15428 6636 16828 6692
rect 16884 6636 16894 6692
rect 17042 6636 17052 6692
rect 17108 6636 18508 6692
rect 18564 6636 18574 6692
rect 21522 6636 21532 6692
rect 21588 6636 22764 6692
rect 22820 6636 22830 6692
rect 22978 6636 22988 6692
rect 23044 6636 24108 6692
rect 24164 6636 24174 6692
rect 24668 6636 25452 6692
rect 25508 6636 27020 6692
rect 27076 6636 33964 6692
rect 34020 6636 34030 6692
rect 38434 6636 38444 6692
rect 38500 6636 39340 6692
rect 39396 6636 39406 6692
rect 22764 6580 22820 6636
rect 4050 6524 4060 6580
rect 4116 6524 4844 6580
rect 4900 6524 5740 6580
rect 5796 6524 5806 6580
rect 5954 6524 5964 6580
rect 6020 6524 6030 6580
rect 8652 6524 9324 6580
rect 9380 6524 16716 6580
rect 16772 6524 16782 6580
rect 17686 6524 17724 6580
rect 17780 6524 17790 6580
rect 22166 6524 22204 6580
rect 22260 6524 22270 6580
rect 22764 6524 25228 6580
rect 25284 6524 25294 6580
rect 27122 6524 27132 6580
rect 27188 6524 29708 6580
rect 29764 6524 30940 6580
rect 30996 6524 31006 6580
rect 31266 6524 31276 6580
rect 31332 6524 32956 6580
rect 33012 6524 33022 6580
rect 39862 6524 39900 6580
rect 39956 6524 42812 6580
rect 42868 6524 42878 6580
rect 4162 6412 4172 6468
rect 4228 6412 5628 6468
rect 5684 6412 6636 6468
rect 6692 6412 6702 6468
rect 8652 6356 8708 6524
rect 30940 6468 30996 6524
rect 8866 6412 8876 6468
rect 8932 6412 9548 6468
rect 9604 6412 10444 6468
rect 10500 6412 18396 6468
rect 18452 6412 18462 6468
rect 20738 6412 20748 6468
rect 20804 6412 20814 6468
rect 22418 6412 22428 6468
rect 22484 6412 23100 6468
rect 23156 6412 23166 6468
rect 23426 6412 23436 6468
rect 23492 6412 25564 6468
rect 25620 6412 25630 6468
rect 27906 6412 27916 6468
rect 27972 6412 28812 6468
rect 28868 6412 28878 6468
rect 30940 6412 35980 6468
rect 36036 6412 36046 6468
rect 38770 6412 38780 6468
rect 38836 6412 41244 6468
rect 41300 6412 41310 6468
rect 20748 6356 20804 6412
rect 3332 6300 8708 6356
rect 16818 6300 16828 6356
rect 16884 6300 17836 6356
rect 17892 6300 17902 6356
rect 20748 6300 22988 6356
rect 23044 6300 26348 6356
rect 26404 6300 26414 6356
rect 29922 6300 29932 6356
rect 29988 6300 33852 6356
rect 33908 6300 33918 6356
rect 36194 6300 36204 6356
rect 36260 6300 41916 6356
rect 41972 6300 41982 6356
rect 3332 6244 3388 6300
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 2706 6188 2716 6244
rect 2772 6188 3388 6244
rect 4610 6188 4620 6244
rect 4676 6188 5404 6244
rect 5460 6188 5470 6244
rect 5618 6188 5628 6244
rect 5684 6188 10332 6244
rect 10388 6188 13468 6244
rect 13524 6188 13534 6244
rect 23762 6188 23772 6244
rect 23828 6188 24220 6244
rect 24276 6188 24286 6244
rect 39554 6188 39564 6244
rect 39620 6188 41804 6244
rect 41860 6188 41870 6244
rect 2034 6076 2044 6132
rect 2100 6076 3164 6132
rect 3220 6076 3230 6132
rect 4946 6076 4956 6132
rect 5012 6076 6748 6132
rect 6804 6076 6814 6132
rect 11554 6076 11564 6132
rect 11620 6076 12124 6132
rect 12180 6076 12190 6132
rect 16818 6076 16828 6132
rect 16884 6076 18284 6132
rect 18340 6076 18350 6132
rect 19506 6076 19516 6132
rect 19572 6076 19852 6132
rect 19908 6076 19918 6132
rect 22642 6076 22652 6132
rect 22708 6076 24444 6132
rect 24500 6076 25564 6132
rect 25620 6076 29036 6132
rect 29092 6076 29102 6132
rect 32722 6076 32732 6132
rect 32788 6076 34412 6132
rect 34468 6076 34478 6132
rect 37202 6076 37212 6132
rect 37268 6076 38220 6132
rect 38276 6076 38286 6132
rect 41682 6076 41692 6132
rect 41748 6076 42140 6132
rect 42196 6076 42206 6132
rect 5394 5964 5404 6020
rect 5460 5964 5516 6020
rect 5572 5964 5582 6020
rect 5730 5964 5740 6020
rect 5796 5964 6972 6020
rect 7028 5964 7038 6020
rect 13570 5964 13580 6020
rect 13636 5964 16156 6020
rect 16212 5964 16222 6020
rect 16902 5964 16940 6020
rect 16996 5964 17006 6020
rect 17602 5964 17612 6020
rect 17668 5964 19068 6020
rect 19124 5964 19134 6020
rect 23958 5964 23996 6020
rect 24052 5964 24062 6020
rect 27346 5964 27356 6020
rect 27412 5964 28476 6020
rect 28532 5964 29260 6020
rect 29316 5964 29326 6020
rect 30940 5964 35084 6020
rect 35140 5964 35150 6020
rect 35970 5964 35980 6020
rect 36036 5964 36876 6020
rect 36932 5964 37772 6020
rect 37828 5964 37838 6020
rect 40086 5964 40124 6020
rect 40180 5964 41132 6020
rect 41188 5964 41198 6020
rect 30940 5908 30996 5964
rect 3938 5852 3948 5908
rect 4004 5852 6524 5908
rect 6580 5852 6590 5908
rect 10210 5852 10220 5908
rect 10276 5852 13356 5908
rect 13412 5852 14476 5908
rect 14532 5852 14542 5908
rect 15026 5852 15036 5908
rect 15092 5852 15820 5908
rect 15876 5852 17948 5908
rect 18004 5852 18014 5908
rect 24434 5852 24444 5908
rect 24500 5852 24892 5908
rect 24948 5852 25788 5908
rect 25844 5852 25854 5908
rect 26310 5852 26348 5908
rect 26404 5852 26414 5908
rect 26674 5852 26684 5908
rect 26740 5852 27580 5908
rect 27636 5852 28364 5908
rect 28420 5852 28430 5908
rect 30930 5852 30940 5908
rect 30996 5852 31006 5908
rect 31490 5852 31500 5908
rect 31556 5852 32396 5908
rect 32452 5852 32462 5908
rect 5170 5740 5180 5796
rect 5236 5740 10164 5796
rect 10322 5740 10332 5796
rect 10388 5740 22204 5796
rect 22260 5740 22270 5796
rect 26114 5740 26124 5796
rect 26180 5740 28252 5796
rect 28308 5740 28318 5796
rect 31042 5740 31052 5796
rect 31108 5740 31724 5796
rect 31780 5740 32060 5796
rect 32116 5740 32126 5796
rect 35746 5740 35756 5796
rect 35812 5740 37436 5796
rect 37492 5740 37502 5796
rect 37762 5740 37772 5796
rect 37828 5740 38892 5796
rect 38948 5740 38958 5796
rect 10108 5684 10164 5740
rect 4834 5628 4844 5684
rect 4900 5628 7308 5684
rect 7364 5628 7374 5684
rect 7858 5628 7868 5684
rect 7924 5628 8428 5684
rect 8484 5628 8494 5684
rect 10108 5628 10556 5684
rect 10612 5628 13468 5684
rect 13524 5628 13534 5684
rect 13906 5628 13916 5684
rect 13972 5628 15372 5684
rect 15428 5628 15438 5684
rect 16930 5628 16940 5684
rect 16996 5628 23660 5684
rect 23716 5628 25340 5684
rect 25396 5628 25406 5684
rect 26852 5628 29372 5684
rect 29428 5628 29438 5684
rect 31826 5628 31836 5684
rect 31892 5628 32620 5684
rect 32676 5628 33180 5684
rect 33236 5628 33246 5684
rect 4022 5516 4060 5572
rect 4116 5516 4126 5572
rect 5282 5516 5292 5572
rect 5348 5516 6300 5572
rect 6356 5516 7980 5572
rect 8036 5516 8316 5572
rect 8372 5516 13692 5572
rect 13748 5516 13758 5572
rect 20300 5516 24220 5572
rect 24276 5516 26572 5572
rect 26628 5516 26638 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 3826 5404 3836 5460
rect 3892 5404 4340 5460
rect 16818 5404 16828 5460
rect 16884 5404 18508 5460
rect 18564 5404 18574 5460
rect 4284 5348 4340 5404
rect 20300 5348 20356 5516
rect 26572 5348 26628 5516
rect 26786 5404 26796 5460
rect 26852 5404 26908 5628
rect 27010 5516 27020 5572
rect 27076 5516 27804 5572
rect 27860 5516 30492 5572
rect 30548 5516 31388 5572
rect 31444 5516 32844 5572
rect 32900 5516 32910 5572
rect 36194 5516 36204 5572
rect 36260 5516 39228 5572
rect 39284 5516 39294 5572
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 27458 5404 27468 5460
rect 27524 5404 28588 5460
rect 28644 5404 31276 5460
rect 31332 5404 32060 5460
rect 32116 5404 32126 5460
rect 35746 5404 35756 5460
rect 35812 5404 35980 5460
rect 36036 5404 39116 5460
rect 39172 5404 39182 5460
rect 3154 5292 3164 5348
rect 3220 5292 3948 5348
rect 4004 5292 4014 5348
rect 4284 5292 4508 5348
rect 4564 5292 4574 5348
rect 12898 5292 12908 5348
rect 12964 5292 20300 5348
rect 20356 5292 20366 5348
rect 24210 5292 24220 5348
rect 24276 5292 26124 5348
rect 26180 5292 26190 5348
rect 26572 5292 28364 5348
rect 28420 5292 29148 5348
rect 29204 5292 29214 5348
rect 35830 5292 35868 5348
rect 35924 5292 37660 5348
rect 37716 5292 37726 5348
rect 38546 5292 38556 5348
rect 38612 5292 41804 5348
rect 41860 5292 41870 5348
rect 2930 5180 2940 5236
rect 2996 5180 5404 5236
rect 5460 5180 5470 5236
rect 6626 5180 6636 5236
rect 6692 5180 8988 5236
rect 9044 5180 9054 5236
rect 15026 5180 15036 5236
rect 15092 5180 15708 5236
rect 15764 5180 15774 5236
rect 17266 5180 17276 5236
rect 17332 5180 18396 5236
rect 18452 5180 18462 5236
rect 20850 5180 20860 5236
rect 20916 5180 21532 5236
rect 21588 5180 21598 5236
rect 23986 5180 23996 5236
rect 24052 5180 25564 5236
rect 25620 5180 25630 5236
rect 25788 5180 27132 5236
rect 27188 5180 27198 5236
rect 28802 5180 28812 5236
rect 28868 5180 31052 5236
rect 31108 5180 32172 5236
rect 32228 5180 32238 5236
rect 32722 5180 32732 5236
rect 32788 5180 33740 5236
rect 33796 5180 33806 5236
rect 36092 5180 37100 5236
rect 37156 5180 37166 5236
rect 41570 5180 41580 5236
rect 41636 5180 41916 5236
rect 41972 5180 41982 5236
rect 25788 5124 25844 5180
rect 36092 5124 36148 5180
rect 3602 5068 3612 5124
rect 3668 5068 5740 5124
rect 5796 5068 5806 5124
rect 12562 5068 12572 5124
rect 12628 5068 13244 5124
rect 13300 5068 19516 5124
rect 19572 5068 21644 5124
rect 21700 5068 21710 5124
rect 25218 5068 25228 5124
rect 25284 5068 25844 5124
rect 26338 5068 26348 5124
rect 26404 5068 27468 5124
rect 27524 5068 27534 5124
rect 34514 5068 34524 5124
rect 34580 5068 36092 5124
rect 36148 5068 36158 5124
rect 36306 5068 36316 5124
rect 36372 5068 36988 5124
rect 37044 5068 37054 5124
rect 41234 5068 41244 5124
rect 41300 5068 41916 5124
rect 41972 5068 41982 5124
rect 26348 5012 26404 5068
rect 4610 4956 4620 5012
rect 4676 4956 7644 5012
rect 7700 4956 7710 5012
rect 11330 4956 11340 5012
rect 11396 4956 12012 5012
rect 12068 4956 12078 5012
rect 12348 4956 14028 5012
rect 14084 4956 14094 5012
rect 18722 4956 18732 5012
rect 18788 4956 19628 5012
rect 19684 4956 19694 5012
rect 23538 4956 23548 5012
rect 23604 4956 24220 5012
rect 24276 4956 24286 5012
rect 24770 4956 24780 5012
rect 24836 4956 26404 5012
rect 26898 4956 26908 5012
rect 26964 4956 30604 5012
rect 30660 4956 30670 5012
rect 30818 4956 30828 5012
rect 30884 4956 32620 5012
rect 32676 4956 32686 5012
rect 39778 4956 39788 5012
rect 39844 4956 41804 5012
rect 41860 4956 41870 5012
rect 4946 4844 4956 4900
rect 5012 4844 7756 4900
rect 7812 4844 7822 4900
rect 10770 4844 10780 4900
rect 10836 4844 12124 4900
rect 12180 4844 12190 4900
rect 12348 4788 12404 4956
rect 4050 4732 4060 4788
rect 4116 4732 6860 4788
rect 6916 4732 6926 4788
rect 8988 4732 10220 4788
rect 10276 4732 10286 4788
rect 11218 4732 11228 4788
rect 11284 4732 12404 4788
rect 13692 4844 15092 4900
rect 23090 4844 23100 4900
rect 23156 4844 24108 4900
rect 24164 4844 24174 4900
rect 39442 4844 39452 4900
rect 39508 4844 40236 4900
rect 40292 4844 40684 4900
rect 40740 4844 40750 4900
rect 8988 4676 9044 4732
rect 13692 4676 13748 4844
rect 1810 4620 1820 4676
rect 1876 4620 9044 4676
rect 9202 4620 9212 4676
rect 9268 4620 13748 4676
rect 15036 4676 15092 4844
rect 22306 4732 22316 4788
rect 22372 4732 23996 4788
rect 24052 4732 24062 4788
rect 37426 4732 37436 4788
rect 37492 4732 38892 4788
rect 38948 4732 42924 4788
rect 42980 4732 42990 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 15036 4620 15484 4676
rect 15540 4620 15596 4676
rect 15652 4620 15662 4676
rect 29026 4620 29036 4676
rect 29092 4620 38332 4676
rect 38388 4620 38398 4676
rect 4722 4508 4732 4564
rect 4788 4508 5404 4564
rect 5460 4508 5470 4564
rect 9090 4508 9100 4564
rect 9156 4508 13860 4564
rect 14018 4508 14028 4564
rect 14084 4508 24724 4564
rect 24882 4508 24892 4564
rect 24948 4508 26012 4564
rect 26068 4508 26078 4564
rect 28130 4508 28140 4564
rect 28196 4508 32844 4564
rect 32900 4508 32910 4564
rect 33394 4508 33404 4564
rect 33460 4508 34972 4564
rect 35028 4508 42252 4564
rect 42308 4508 42318 4564
rect 13804 4452 13860 4508
rect 24668 4452 24724 4508
rect 3938 4396 3948 4452
rect 4004 4396 5852 4452
rect 5908 4396 5918 4452
rect 11106 4396 11116 4452
rect 11172 4396 11900 4452
rect 11956 4396 11966 4452
rect 12674 4396 12684 4452
rect 12740 4396 13580 4452
rect 13636 4396 13646 4452
rect 13804 4396 18732 4452
rect 18788 4396 18798 4452
rect 24668 4396 25452 4452
rect 25508 4396 26572 4452
rect 26628 4396 26638 4452
rect 30034 4396 30044 4452
rect 30100 4396 30716 4452
rect 30772 4396 30782 4452
rect 38770 4396 38780 4452
rect 38836 4396 40124 4452
rect 40180 4396 40190 4452
rect 3714 4284 3724 4340
rect 3780 4284 17164 4340
rect 17220 4284 17230 4340
rect 24098 4284 24108 4340
rect 24164 4284 26460 4340
rect 26516 4284 29932 4340
rect 29988 4284 32284 4340
rect 32340 4284 36428 4340
rect 36484 4284 36494 4340
rect 36652 4284 41580 4340
rect 41636 4284 41804 4340
rect 41860 4284 41870 4340
rect 36652 4228 36708 4284
rect 1138 4172 1148 4228
rect 1204 4172 1932 4228
rect 1988 4172 1998 4228
rect 5170 4172 5180 4228
rect 5236 4172 6076 4228
rect 6132 4172 6142 4228
rect 7298 4172 7308 4228
rect 7364 4172 12908 4228
rect 12964 4172 12974 4228
rect 14578 4172 14588 4228
rect 14644 4172 15484 4228
rect 15540 4172 15550 4228
rect 21298 4172 21308 4228
rect 21364 4172 21374 4228
rect 22194 4172 22204 4228
rect 22260 4172 24892 4228
rect 24948 4172 24958 4228
rect 31826 4172 31836 4228
rect 31892 4172 33628 4228
rect 33684 4172 36708 4228
rect 38612 4172 39676 4228
rect 39732 4172 39742 4228
rect 7308 4116 7364 4172
rect 21308 4116 21364 4172
rect 38612 4116 38668 4172
rect 3826 4060 3836 4116
rect 3892 4060 5964 4116
rect 6020 4060 7364 4116
rect 13234 4060 13244 4116
rect 13300 4060 21364 4116
rect 34290 4060 34300 4116
rect 34356 4060 35532 4116
rect 35588 4060 38668 4116
rect 21298 3948 21308 4004
rect 21364 3948 22316 4004
rect 22372 3948 22382 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23986 3724 23996 3780
rect 24052 3724 26348 3780
rect 26404 3724 26414 3780
rect 34514 3724 34524 3780
rect 34580 3724 35756 3780
rect 35812 3724 37772 3780
rect 37828 3724 37838 3780
rect 38612 3724 39004 3780
rect 39060 3724 39070 3780
rect 39778 3724 39788 3780
rect 39844 3724 41580 3780
rect 41636 3724 42364 3780
rect 42420 3724 42430 3780
rect 38612 3668 38668 3724
rect 13234 3612 13244 3668
rect 13300 3612 14252 3668
rect 14308 3612 14318 3668
rect 17826 3612 17836 3668
rect 17892 3612 21532 3668
rect 21588 3612 21598 3668
rect 24210 3612 24220 3668
rect 24276 3612 29260 3668
rect 29316 3612 29326 3668
rect 31378 3612 31388 3668
rect 31444 3612 35868 3668
rect 35924 3612 38668 3668
rect 4834 3500 4844 3556
rect 4900 3500 9772 3556
rect 9828 3500 9838 3556
rect 14130 3500 14140 3556
rect 14196 3500 17612 3556
rect 17668 3500 17678 3556
rect 23426 3500 23436 3556
rect 23492 3500 26068 3556
rect 26898 3500 26908 3556
rect 26964 3500 27580 3556
rect 27636 3500 27646 3556
rect 38322 3500 38332 3556
rect 38388 3500 39116 3556
rect 39172 3500 39182 3556
rect 39554 3500 39564 3556
rect 39620 3500 40908 3556
rect 40964 3500 40974 3556
rect 41346 3500 41356 3556
rect 41412 3500 41468 3556
rect 41524 3500 41534 3556
rect 26012 3444 26068 3500
rect 41356 3444 41412 3500
rect 24994 3388 25004 3444
rect 25060 3388 25788 3444
rect 25844 3388 25854 3444
rect 26012 3388 26684 3444
rect 26740 3388 30268 3444
rect 30324 3388 30334 3444
rect 34738 3388 34748 3444
rect 34804 3388 38108 3444
rect 38164 3388 38174 3444
rect 39330 3388 39340 3444
rect 39396 3388 41412 3444
rect 4162 3276 4172 3332
rect 4228 3276 25004 3332
rect 25060 3276 25070 3332
rect 32498 3276 32508 3332
rect 32564 3276 37212 3332
rect 37268 3276 37278 3332
rect 38612 3276 40124 3332
rect 40180 3276 40190 3332
rect 41458 3276 41468 3332
rect 41524 3276 41534 3332
rect 38612 3220 38668 3276
rect 35410 3164 35420 3220
rect 35476 3164 38668 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 41468 3108 41524 3276
rect 22082 3052 22092 3108
rect 22148 3052 23044 3108
rect 36530 3052 36540 3108
rect 36596 3052 41524 3108
rect 22988 2996 23044 3052
rect 3490 2940 3500 2996
rect 3556 2940 22652 2996
rect 22708 2940 22718 2996
rect 22988 2940 38780 2996
rect 38836 2940 38846 2996
rect 24658 2828 24668 2884
rect 24724 2828 35420 2884
rect 35476 2828 35486 2884
rect 38434 2828 38444 2884
rect 38500 2828 43036 2884
rect 43092 2828 43102 2884
rect 24882 2716 24892 2772
rect 24948 2716 37324 2772
rect 37380 2716 37390 2772
rect 1586 2604 1596 2660
rect 1652 2604 29372 2660
rect 29428 2604 29438 2660
rect 35298 2604 35308 2660
rect 35364 2604 43372 2660
rect 43428 2604 43438 2660
rect 31154 2492 31164 2548
rect 31220 2492 42588 2548
rect 42644 2492 42654 2548
rect 1698 2380 1708 2436
rect 1764 2380 34748 2436
rect 34804 2380 34814 2436
rect 36082 2044 36092 2100
rect 36148 2044 38444 2100
rect 38500 2044 38510 2100
rect 25778 1596 25788 1652
rect 25844 1596 38668 1652
rect 38724 1596 38734 1652
rect 32050 1484 32060 1540
rect 32116 1484 34524 1540
rect 34580 1484 42700 1540
rect 42756 1484 42766 1540
<< via3 >>
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 18396 23996 18452 24052
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 32620 23660 32676 23716
rect 39340 23660 39396 23716
rect 40124 23660 40180 23716
rect 39900 23548 39956 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 40012 22988 40068 23044
rect 28812 22876 28868 22932
rect 30604 22876 30660 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 29484 22316 29540 22372
rect 40684 22204 40740 22260
rect 30604 22092 30660 22148
rect 34972 22092 35028 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 29372 21868 29428 21924
rect 40684 21868 40740 21924
rect 28924 21756 28980 21812
rect 33516 21644 33572 21700
rect 23436 21420 23492 21476
rect 25564 21420 25620 21476
rect 30716 21420 30772 21476
rect 25116 21308 25172 21364
rect 33740 21308 33796 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 34748 21084 34804 21140
rect 32732 20860 32788 20916
rect 26684 20748 26740 20804
rect 36092 20748 36148 20804
rect 29148 20636 29204 20692
rect 32732 20636 32788 20692
rect 33516 20636 33572 20692
rect 30268 20524 30324 20580
rect 34300 20524 34356 20580
rect 34748 20524 34804 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 33292 20300 33348 20356
rect 36316 20300 36372 20356
rect 39676 20300 39732 20356
rect 26124 20076 26180 20132
rect 28364 20076 28420 20132
rect 33292 20076 33348 20132
rect 22092 19852 22148 19908
rect 24668 19852 24724 19908
rect 27356 19852 27412 19908
rect 34972 19852 35028 19908
rect 36764 19852 36820 19908
rect 38444 19852 38500 19908
rect 27132 19740 27188 19796
rect 30940 19740 30996 19796
rect 36316 19740 36372 19796
rect 36988 19628 37044 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 33852 19404 33908 19460
rect 34524 19292 34580 19348
rect 36428 19180 36484 19236
rect 27356 19068 27412 19124
rect 22204 18956 22260 19012
rect 37436 18844 37492 18900
rect 38892 18844 38948 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 28476 18508 28532 18564
rect 31164 18508 31220 18564
rect 35868 18508 35924 18564
rect 31612 18284 31668 18340
rect 34972 18172 35028 18228
rect 36428 18172 36484 18228
rect 41356 18172 41412 18228
rect 41244 18060 41300 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 29820 17948 29876 18004
rect 30268 17948 30324 18004
rect 37212 17948 37268 18004
rect 42364 17948 42420 18004
rect 34412 17836 34468 17892
rect 31276 17724 31332 17780
rect 41916 17724 41972 17780
rect 27356 17388 27412 17444
rect 38332 17388 38388 17444
rect 41356 17388 41412 17444
rect 25564 17276 25620 17332
rect 33964 17276 34020 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 27580 16940 27636 16996
rect 15484 16828 15540 16884
rect 16940 16828 16996 16884
rect 25564 16828 25620 16884
rect 26348 16828 26404 16884
rect 29036 16828 29092 16884
rect 33628 17164 33684 17220
rect 41244 17052 41300 17108
rect 39116 16940 39172 16996
rect 39228 16604 39284 16660
rect 33292 16492 33348 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 28252 16380 28308 16436
rect 41916 16380 41972 16436
rect 25116 16268 25172 16324
rect 41468 16268 41524 16324
rect 31164 16156 31220 16212
rect 39116 16044 39172 16100
rect 27356 15932 27412 15988
rect 28252 15932 28308 15988
rect 34860 15932 34916 15988
rect 40572 15932 40628 15988
rect 41692 15820 41748 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 32172 15596 32228 15652
rect 38220 15596 38276 15652
rect 39452 15484 39508 15540
rect 38444 15260 38500 15316
rect 35868 15148 35924 15204
rect 32172 14924 32228 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 28476 14812 28532 14868
rect 38668 14812 38724 14868
rect 33852 14700 33908 14756
rect 31388 14588 31444 14644
rect 27132 14476 27188 14532
rect 41916 14476 41972 14532
rect 36652 14252 36708 14308
rect 31388 14140 31444 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 33852 14140 33908 14196
rect 42364 14028 42420 14084
rect 28364 13916 28420 13972
rect 39564 13916 39620 13972
rect 41692 13916 41748 13972
rect 30492 13692 30548 13748
rect 33292 13692 33348 13748
rect 36764 13692 36820 13748
rect 38220 13692 38276 13748
rect 34972 13580 35028 13636
rect 38108 13580 38164 13636
rect 13916 13468 13972 13524
rect 24668 13356 24724 13412
rect 30828 13356 30884 13412
rect 32284 13356 32340 13412
rect 34860 13356 34916 13412
rect 40572 13356 40628 13412
rect 41580 13356 41636 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 29148 13244 29204 13300
rect 38780 13132 38836 13188
rect 40012 13132 40068 13188
rect 30828 13020 30884 13076
rect 32844 12908 32900 12964
rect 36988 12908 37044 12964
rect 41468 12908 41524 12964
rect 31612 12796 31668 12852
rect 34300 12796 34356 12852
rect 30940 12684 30996 12740
rect 33740 12684 33796 12740
rect 34748 12684 34804 12740
rect 26908 12572 26964 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 30716 12460 30772 12516
rect 31052 12460 31108 12516
rect 12796 12348 12852 12404
rect 10332 12236 10388 12292
rect 29820 12348 29876 12404
rect 31388 12348 31444 12404
rect 33516 12348 33572 12404
rect 38332 12348 38388 12404
rect 39564 12348 39620 12404
rect 17052 12236 17108 12292
rect 27580 12236 27636 12292
rect 34300 12236 34356 12292
rect 34524 12236 34580 12292
rect 36988 12236 37044 12292
rect 13468 12124 13524 12180
rect 16828 12124 16884 12180
rect 29148 12124 29204 12180
rect 31164 12124 31220 12180
rect 30492 12012 30548 12068
rect 30828 12012 30884 12068
rect 31052 12012 31108 12068
rect 33964 12012 34020 12068
rect 34300 12012 34356 12068
rect 37436 12012 37492 12068
rect 31164 11900 31220 11956
rect 32284 11788 32340 11844
rect 38668 11788 38724 11844
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 31164 11732 31220 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 12796 11676 12852 11732
rect 37324 11676 37380 11732
rect 16604 11564 16660 11620
rect 17052 11564 17108 11620
rect 26908 11564 26964 11620
rect 35756 11564 35812 11620
rect 38892 11564 38948 11620
rect 13916 11452 13972 11508
rect 28924 11452 28980 11508
rect 32844 11340 32900 11396
rect 39788 11340 39844 11396
rect 18396 11228 18452 11284
rect 34300 11228 34356 11284
rect 34636 11228 34692 11284
rect 37212 11228 37268 11284
rect 37436 11116 37492 11172
rect 37660 11116 37716 11172
rect 38892 11116 38948 11172
rect 41692 11116 41748 11172
rect 39788 11004 39844 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 13916 10892 13972 10948
rect 17724 10892 17780 10948
rect 19516 10892 19572 10948
rect 35980 10892 36036 10948
rect 24668 10780 24724 10836
rect 34636 10780 34692 10836
rect 36428 10780 36484 10836
rect 17500 10444 17556 10500
rect 36652 10332 36708 10388
rect 39340 10332 39396 10388
rect 17612 10220 17668 10276
rect 37436 10220 37492 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 16604 10108 16660 10164
rect 32844 10108 32900 10164
rect 34300 10108 34356 10164
rect 34636 10108 34692 10164
rect 38220 10108 38276 10164
rect 17500 9996 17556 10052
rect 22316 9996 22372 10052
rect 29484 9884 29540 9940
rect 35644 9884 35700 9940
rect 36092 9772 36148 9828
rect 40684 9772 40740 9828
rect 37436 9660 37492 9716
rect 41580 9660 41636 9716
rect 16828 9548 16884 9604
rect 26684 9548 26740 9604
rect 38780 9548 38836 9604
rect 39788 9548 39844 9604
rect 26460 9436 26516 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 39564 9436 39620 9492
rect 17612 9324 17668 9380
rect 35868 9324 35924 9380
rect 5292 9212 5348 9268
rect 17052 9212 17108 9268
rect 29036 9212 29092 9268
rect 39676 9212 39732 9268
rect 41916 9212 41972 9268
rect 26124 9100 26180 9156
rect 26460 9100 26516 9156
rect 36428 9100 36484 9156
rect 5180 8988 5236 9044
rect 34748 8988 34804 9044
rect 38220 8988 38276 9044
rect 39788 8876 39844 8932
rect 37324 8764 37380 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 24668 8540 24724 8596
rect 36428 8540 36484 8596
rect 10332 8428 10388 8484
rect 5404 8316 5460 8372
rect 29372 8316 29428 8372
rect 36316 8204 36372 8260
rect 38108 8204 38164 8260
rect 29372 8092 29428 8148
rect 41692 8092 41748 8148
rect 5852 7980 5908 8036
rect 30604 7980 30660 8036
rect 36316 7868 36372 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 33628 7756 33684 7812
rect 35644 7756 35700 7812
rect 30716 7644 30772 7700
rect 5180 7308 5236 7364
rect 34636 7308 34692 7364
rect 5628 7196 5684 7252
rect 28812 7196 28868 7252
rect 30716 7196 30772 7252
rect 5292 7084 5348 7140
rect 23996 7084 24052 7140
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 16604 6972 16660 7028
rect 13468 6860 13524 6916
rect 39340 6636 39396 6692
rect 4060 6524 4116 6580
rect 5740 6524 5796 6580
rect 17724 6524 17780 6580
rect 22204 6524 22260 6580
rect 39900 6524 39956 6580
rect 28812 6412 28868 6468
rect 33852 6300 33908 6356
rect 41916 6300 41972 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 5404 6188 5460 6244
rect 5628 6188 5684 6244
rect 13468 6188 13524 6244
rect 39564 6188 39620 6244
rect 19516 6076 19572 6132
rect 34412 6076 34468 6132
rect 5404 5964 5460 6020
rect 16940 5964 16996 6020
rect 23996 5964 24052 6020
rect 40124 5964 40180 6020
rect 26348 5852 26404 5908
rect 16940 5628 16996 5684
rect 4060 5516 4116 5572
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 39228 5516 39284 5572
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 35980 5404 36036 5460
rect 35868 5292 35924 5348
rect 41916 5180 41972 5236
rect 26348 5068 26404 5124
rect 30604 4956 30660 5012
rect 32620 4956 32676 5012
rect 39452 4844 39508 4900
rect 22316 4732 22372 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 15484 4620 15540 4676
rect 5404 4508 5460 4564
rect 41580 4284 41636 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 34524 3724 34580 3780
rect 31388 3612 31444 3668
rect 23436 3500 23492 3556
rect 41468 3500 41524 3556
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 22092 3052 22148 3108
rect 37324 2716 37380 2772
<< metal4 >>
rect 4448 40012 4768 40828
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 19808 40796 20128 40828
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 18396 24052 18452 24062
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 15484 16884 15540 16894
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 13916 13524 13972 13534
rect 12796 12404 12852 12414
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 10332 12292 10388 12302
rect 5292 9268 5348 9278
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 5180 9044 5236 9054
rect 5180 7364 5236 8988
rect 5180 7298 5236 7308
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 5292 7140 5348 9212
rect 10332 8484 10388 12236
rect 12796 11732 12852 12348
rect 12796 11666 12852 11676
rect 13468 12180 13524 12190
rect 10332 8418 10388 8428
rect 5292 7074 5348 7084
rect 5404 8372 5460 8382
rect 4060 6580 4116 6590
rect 4060 5572 4116 6524
rect 4060 5506 4116 5516
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 5404 6244 5460 8316
rect 5852 8036 5908 8046
rect 5740 7980 5852 8036
rect 5404 6020 5460 6188
rect 5628 7252 5684 7262
rect 5628 6244 5684 7196
rect 5740 6580 5796 7980
rect 5852 7970 5908 7980
rect 5740 6514 5796 6524
rect 13468 6916 13524 12124
rect 13916 11508 13972 13468
rect 13916 10948 13972 11452
rect 13916 10882 13972 10892
rect 5628 6178 5684 6188
rect 13468 6244 13524 6860
rect 13468 6178 13524 6188
rect 5404 4564 5460 5964
rect 15484 4676 15540 16828
rect 16940 16884 16996 16894
rect 16828 12180 16884 12190
rect 16604 11620 16660 11630
rect 16604 10164 16660 11564
rect 16604 7028 16660 10108
rect 16828 9604 16884 12124
rect 16828 9538 16884 9548
rect 16604 6962 16660 6972
rect 16940 6020 16996 16828
rect 17052 12292 17108 12302
rect 17052 11620 17108 12236
rect 17052 9268 17108 11564
rect 18396 11284 18452 23996
rect 18396 11218 18452 11228
rect 19808 23548 20128 25060
rect 35168 40012 35488 40828
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 32620 23716 32676 23726
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 28812 22932 28868 22942
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 23436 21476 23492 21486
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 17724 10948 17780 10958
rect 17500 10500 17556 10510
rect 17500 10052 17556 10444
rect 17500 9986 17556 9996
rect 17612 10276 17668 10286
rect 17612 9380 17668 10220
rect 17612 9314 17668 9324
rect 17052 9202 17108 9212
rect 17724 6580 17780 10892
rect 17724 6514 17780 6524
rect 19516 10948 19572 10958
rect 19516 6132 19572 10892
rect 19516 6066 19572 6076
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 16940 5684 16996 5964
rect 16940 5618 16996 5628
rect 15484 4610 15540 4620
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 5404 4498 5460 4508
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 22092 19908 22148 19918
rect 22092 3108 22148 19852
rect 22204 19012 22260 19022
rect 22204 6580 22260 18956
rect 22204 6514 22260 6524
rect 22316 10052 22372 10062
rect 22316 4788 22372 9996
rect 22316 4722 22372 4732
rect 23436 3556 23492 21420
rect 25564 21476 25620 21486
rect 25116 21364 25172 21374
rect 24668 19908 24724 19918
rect 24668 13412 24724 19852
rect 25116 16324 25172 21308
rect 25564 17332 25620 21420
rect 26684 20804 26740 20814
rect 25564 16884 25620 17276
rect 25564 16818 25620 16828
rect 26124 20132 26180 20142
rect 25116 16258 25172 16268
rect 24668 13346 24724 13356
rect 24668 10836 24724 10846
rect 24668 8596 24724 10780
rect 26124 9156 26180 20076
rect 26124 9090 26180 9100
rect 26348 16884 26404 16894
rect 24668 8530 24724 8540
rect 23996 7140 24052 7150
rect 23996 6020 24052 7084
rect 23996 5954 24052 5964
rect 26348 5908 26404 16828
rect 26684 9604 26740 20748
rect 28364 20132 28420 20142
rect 27356 19908 27412 19918
rect 27132 19796 27188 19806
rect 27132 14532 27188 19740
rect 27356 19124 27412 19852
rect 27356 19058 27412 19068
rect 27356 17444 27412 17454
rect 27356 15988 27412 17388
rect 27356 15922 27412 15932
rect 27580 16996 27636 17006
rect 27132 14466 27188 14476
rect 26908 12628 26964 12638
rect 26908 11620 26964 12572
rect 27580 12292 27636 16940
rect 28252 16436 28308 16446
rect 28252 15988 28308 16380
rect 28252 15922 28308 15932
rect 28364 13972 28420 20076
rect 28476 18564 28532 18574
rect 28476 14868 28532 18508
rect 28476 14802 28532 14812
rect 28364 13906 28420 13916
rect 27580 12226 27636 12236
rect 26908 11554 26964 11564
rect 26684 9538 26740 9548
rect 26460 9492 26516 9502
rect 26460 9156 26516 9436
rect 26460 9090 26516 9100
rect 28812 7252 28868 22876
rect 30604 22932 30660 22942
rect 29484 22372 29540 22382
rect 29372 21924 29428 21934
rect 28924 21812 28980 21822
rect 28924 11508 28980 21756
rect 29148 20692 29204 20702
rect 28924 11442 28980 11452
rect 29036 16884 29092 16894
rect 29036 9268 29092 16828
rect 29148 13300 29204 20636
rect 29148 12180 29204 13244
rect 29148 12114 29204 12124
rect 29036 9202 29092 9212
rect 29372 8372 29428 21868
rect 29484 9940 29540 22316
rect 30604 22148 30660 22876
rect 30268 20580 30324 20590
rect 29820 18004 29876 18014
rect 29820 12404 29876 17948
rect 30268 18004 30324 20524
rect 30268 17938 30324 17948
rect 29820 12338 29876 12348
rect 30492 13748 30548 13758
rect 30492 12068 30548 13692
rect 30492 12002 30548 12012
rect 29484 9874 29540 9884
rect 29372 8148 29428 8316
rect 29372 8082 29428 8092
rect 28812 6468 28868 7196
rect 28812 6402 28868 6412
rect 30604 8036 30660 22092
rect 30716 21476 30772 21486
rect 30716 12516 30772 21420
rect 30940 19796 30996 19806
rect 30828 13412 30884 13422
rect 30828 13076 30884 13356
rect 30828 13010 30884 13020
rect 30940 12740 30996 19740
rect 30716 12450 30772 12460
rect 30828 12684 30940 12740
rect 30828 12068 30884 12684
rect 30940 12674 30996 12684
rect 31164 18564 31220 18574
rect 31164 16212 31220 18508
rect 31612 18340 31668 18350
rect 30828 12002 30884 12012
rect 31052 12516 31108 12526
rect 31052 12068 31108 12460
rect 31164 12180 31220 16156
rect 31276 17780 31332 17790
rect 31276 15148 31332 17724
rect 31276 15092 31444 15148
rect 31388 14644 31444 15092
rect 31388 14196 31444 14588
rect 31388 14130 31444 14140
rect 31612 12852 31668 18284
rect 32172 15652 32228 15662
rect 32172 14980 32228 15596
rect 32172 14914 32228 14924
rect 31612 12786 31668 12796
rect 32284 13412 32340 13422
rect 31164 12114 31220 12124
rect 31388 12404 31444 12414
rect 31052 12002 31108 12012
rect 31164 11956 31220 11966
rect 31164 11788 31220 11900
rect 31164 11722 31220 11732
rect 26348 5124 26404 5852
rect 26348 5058 26404 5068
rect 30604 5012 30660 7980
rect 30716 7700 30772 7710
rect 30716 7252 30772 7644
rect 30716 7186 30772 7196
rect 30604 4946 30660 4956
rect 31388 3668 31444 12348
rect 32284 11844 32340 13356
rect 32284 11778 32340 11788
rect 32620 5012 32676 23660
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 34972 22148 35028 22158
rect 33516 21700 33572 21710
rect 32732 20916 32788 20926
rect 32732 20692 32788 20860
rect 32732 20626 32788 20636
rect 33516 20692 33572 21644
rect 33292 20356 33348 20366
rect 33292 20132 33348 20300
rect 33292 20066 33348 20076
rect 33292 16548 33348 16558
rect 33292 13748 33348 16492
rect 33292 13682 33348 13692
rect 32844 12964 32900 12974
rect 32844 11396 32900 12908
rect 33516 12404 33572 20636
rect 33740 21364 33796 21374
rect 33516 12338 33572 12348
rect 33628 17220 33684 17230
rect 32844 10164 32900 11340
rect 32844 10098 32900 10108
rect 33628 7812 33684 17164
rect 33740 12740 33796 21308
rect 34748 21140 34804 21150
rect 34300 20580 34356 20590
rect 33852 19460 33908 19470
rect 33852 14756 33908 19404
rect 33852 14690 33908 14700
rect 33964 17332 34020 17342
rect 33740 12674 33796 12684
rect 33852 14196 33908 14206
rect 33628 7746 33684 7756
rect 33852 6356 33908 14140
rect 33964 12068 34020 17276
rect 33964 12002 34020 12012
rect 34300 12852 34356 20524
rect 34748 20580 34804 21084
rect 34524 19348 34580 19358
rect 34300 12292 34356 12796
rect 34300 12068 34356 12236
rect 34300 12002 34356 12012
rect 34412 17892 34468 17902
rect 34300 11284 34356 11294
rect 34300 10164 34356 11228
rect 34300 10098 34356 10108
rect 33852 6290 33908 6300
rect 34412 6132 34468 17836
rect 34412 6066 34468 6076
rect 34524 12292 34580 19292
rect 34748 15148 34804 20524
rect 34972 19908 35028 22092
rect 34972 19842 35028 19852
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 39340 23716 39396 23726
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 34972 18228 35028 18238
rect 32620 4946 32676 4956
rect 34524 3780 34580 12236
rect 34636 15092 34804 15148
rect 34860 15988 34916 15998
rect 34636 11284 34692 15092
rect 34860 13412 34916 15932
rect 34972 13636 35028 18172
rect 34972 13570 35028 13580
rect 35168 18060 35488 19572
rect 36092 20804 36148 20814
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35868 18564 35924 18574
rect 35868 15204 35924 18508
rect 35868 15138 35924 15148
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 34860 13346 34916 13356
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 34636 11218 34692 11228
rect 34748 12740 34804 12750
rect 34636 10836 34692 10846
rect 34636 10164 34692 10780
rect 34636 7364 34692 10108
rect 34748 9044 34804 12684
rect 34748 8978 34804 8988
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 34636 7298 34692 7308
rect 35168 8652 35488 10164
rect 35756 11620 35812 11630
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 34524 3714 34580 3724
rect 35168 7084 35488 8596
rect 35644 9940 35700 9950
rect 35756 9940 35812 11564
rect 35700 9884 35812 9940
rect 35980 10948 36036 10958
rect 35644 7812 35700 9884
rect 35644 7746 35700 7756
rect 35868 9380 35924 9390
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35868 5348 35924 9324
rect 35980 5460 36036 10892
rect 36092 9828 36148 20748
rect 36316 20356 36372 20366
rect 36316 19796 36372 20300
rect 36316 19730 36372 19740
rect 36764 19908 36820 19918
rect 36428 19236 36484 19246
rect 36428 18228 36484 19180
rect 36428 10836 36484 18172
rect 36428 10770 36484 10780
rect 36652 14308 36708 14318
rect 36652 10388 36708 14252
rect 36764 13748 36820 19852
rect 38444 19908 38500 19918
rect 36764 13682 36820 13692
rect 36988 19684 37044 19694
rect 36988 12964 37044 19628
rect 37436 18900 37492 18910
rect 36988 12292 37044 12908
rect 36988 12226 37044 12236
rect 37212 18004 37268 18014
rect 37212 11284 37268 17948
rect 37436 12068 37492 18844
rect 38332 17444 38388 17454
rect 38220 15652 38276 15662
rect 38220 13748 38276 15596
rect 38220 13682 38276 13692
rect 37436 12002 37492 12012
rect 38108 13636 38164 13646
rect 37324 11732 37380 11742
rect 37380 11676 37716 11732
rect 37324 11666 37380 11676
rect 37212 11218 37268 11228
rect 36652 10322 36708 10332
rect 37436 11172 37492 11182
rect 36092 9762 36148 9772
rect 37436 10276 37492 11116
rect 37660 11172 37716 11676
rect 37660 11106 37716 11116
rect 37436 9716 37492 10220
rect 37436 9650 37492 9660
rect 36428 9156 36484 9166
rect 36428 8596 36484 9100
rect 36428 8530 36484 8540
rect 37324 8820 37380 8830
rect 36316 8260 36372 8270
rect 36316 7924 36372 8204
rect 36316 7858 36372 7868
rect 35980 5394 36036 5404
rect 35868 5282 35924 5292
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 31388 3602 31444 3612
rect 23436 3490 23492 3500
rect 35168 3076 35488 3892
rect 22092 3042 22148 3052
rect 37324 2772 37380 8764
rect 38108 8260 38164 13580
rect 38332 12404 38388 17388
rect 38444 15316 38500 19852
rect 38444 15250 38500 15260
rect 38892 18900 38948 18910
rect 38332 12338 38388 12348
rect 38668 14868 38724 14878
rect 38668 11844 38724 14812
rect 38668 11778 38724 11788
rect 38780 13188 38836 13198
rect 38220 10164 38276 10174
rect 38220 9044 38276 10108
rect 38780 9604 38836 13132
rect 38892 11620 38948 18844
rect 39116 16996 39172 17006
rect 39116 16100 39172 16940
rect 39116 16034 39172 16044
rect 39228 16660 39284 16670
rect 38892 11172 38948 11564
rect 38892 11106 38948 11116
rect 38780 9538 38836 9548
rect 38220 8978 38276 8988
rect 38108 8194 38164 8204
rect 39228 5572 39284 16604
rect 39340 10612 39396 23660
rect 40124 23716 40180 23726
rect 39900 23604 39956 23614
rect 39676 20356 39732 20366
rect 39452 15540 39508 15550
rect 39452 11788 39508 15484
rect 39564 13972 39620 13982
rect 39564 12404 39620 13916
rect 39564 12338 39620 12348
rect 39452 11732 39620 11788
rect 39340 10556 39508 10612
rect 39340 10388 39396 10398
rect 39340 6692 39396 10332
rect 39340 6626 39396 6636
rect 39228 5506 39284 5516
rect 39452 4900 39508 10556
rect 39564 9492 39620 11732
rect 39564 6244 39620 9436
rect 39676 9268 39732 20300
rect 39788 11396 39844 11406
rect 39788 11060 39844 11340
rect 39788 10994 39844 11004
rect 39676 9202 39732 9212
rect 39788 9604 39844 9614
rect 39788 8932 39844 9548
rect 39788 8866 39844 8876
rect 39900 6580 39956 23548
rect 40012 23044 40068 23054
rect 40012 13188 40068 22988
rect 40012 13122 40068 13132
rect 39900 6514 39956 6524
rect 39564 6178 39620 6188
rect 40124 6020 40180 23660
rect 40684 22260 40740 22270
rect 40684 21924 40740 22204
rect 40572 15988 40628 15998
rect 40572 13412 40628 15932
rect 40572 13346 40628 13356
rect 40684 9828 40740 21868
rect 41356 18228 41412 18238
rect 41244 18116 41300 18126
rect 41244 17108 41300 18060
rect 41356 17444 41412 18172
rect 42364 18004 42420 18014
rect 41356 17378 41412 17388
rect 41916 17780 41972 17790
rect 41244 17042 41300 17052
rect 41916 16436 41972 17724
rect 41916 16370 41972 16380
rect 40684 9762 40740 9772
rect 41468 16324 41524 16334
rect 41468 12964 41524 16268
rect 41692 15876 41748 15886
rect 41692 13972 41748 15820
rect 41692 13906 41748 13916
rect 41916 14532 41972 14542
rect 40124 5954 40180 5964
rect 39452 4834 39508 4844
rect 41468 3556 41524 12908
rect 41580 13412 41636 13422
rect 41580 9716 41636 13356
rect 41580 4340 41636 9660
rect 41692 11172 41748 11182
rect 41692 8148 41748 11116
rect 41692 8082 41748 8092
rect 41916 9268 41972 14476
rect 42364 14084 42420 17948
rect 42364 14018 42420 14028
rect 41916 6356 41972 9212
rect 41916 5236 41972 6300
rect 41916 5170 41972 5180
rect 41580 4274 41636 4284
rect 41468 3490 41524 3500
rect 37324 2706 37380 2716
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__I gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A1
timestamp 1669390400
transform 1 0 29904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__A2
timestamp 1669390400
transform 1 0 30464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__I
timestamp 1669390400
transform 1 0 15568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__I
timestamp 1669390400
transform -1 0 14000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__A1
timestamp 1669390400
transform 1 0 4032 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__A2
timestamp 1669390400
transform 1 0 5936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__I
timestamp 1669390400
transform -1 0 37296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A1
timestamp 1669390400
transform -1 0 2800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__A1
timestamp 1669390400
transform 1 0 5040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__A1
timestamp 1669390400
transform -1 0 3248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__I
timestamp 1669390400
transform 1 0 33488 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A1
timestamp 1669390400
transform 1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__A2
timestamp 1669390400
transform -1 0 4816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A1
timestamp 1669390400
transform -1 0 2240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__A2
timestamp 1669390400
transform -1 0 2912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1669390400
transform 1 0 3360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__I
timestamp 1669390400
transform 1 0 11424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A1
timestamp 1669390400
transform 1 0 3584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__A2
timestamp 1669390400
transform -1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__I
timestamp 1669390400
transform -1 0 4144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__A1
timestamp 1669390400
transform 1 0 5600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__371__I
timestamp 1669390400
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__A1
timestamp 1669390400
transform 1 0 13328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__372__A2
timestamp 1669390400
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A1
timestamp 1669390400
transform 1 0 15680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__373__A2
timestamp 1669390400
transform -1 0 3920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__375__I
timestamp 1669390400
transform 1 0 17360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A1
timestamp 1669390400
transform 1 0 4480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A2
timestamp 1669390400
transform 1 0 2800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A1
timestamp 1669390400
transform 1 0 14560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__A2
timestamp 1669390400
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__380__A1
timestamp 1669390400
transform 1 0 14336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__382__A1
timestamp 1669390400
transform 1 0 17808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__384__A1
timestamp 1669390400
transform 1 0 16016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A1
timestamp 1669390400
transform 1 0 37968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2
timestamp 1669390400
transform 1 0 38752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1669390400
transform -1 0 10416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A1
timestamp 1669390400
transform 1 0 19936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__388__A2
timestamp 1669390400
transform 1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__389__I
timestamp 1669390400
transform 1 0 28224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__I
timestamp 1669390400
transform -1 0 17360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A1
timestamp 1669390400
transform -1 0 19152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__A2
timestamp 1669390400
transform -1 0 16912 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__391__B
timestamp 1669390400
transform 1 0 20832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A1
timestamp 1669390400
transform -1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__392__A2
timestamp 1669390400
transform 1 0 19040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__393__A4
timestamp 1669390400
transform -1 0 36512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A1
timestamp 1669390400
transform -1 0 41328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__395__A2
timestamp 1669390400
transform -1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A1
timestamp 1669390400
transform -1 0 25312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A2
timestamp 1669390400
transform -1 0 23520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A3
timestamp 1669390400
transform -1 0 22624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__396__A4
timestamp 1669390400
transform -1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__397__A1
timestamp 1669390400
transform -1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1
timestamp 1669390400
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1669390400
transform -1 0 9856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A3
timestamp 1669390400
transform -1 0 25312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A1
timestamp 1669390400
transform 1 0 15792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__399__A2
timestamp 1669390400
transform 1 0 16240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__400__A2
timestamp 1669390400
transform 1 0 17584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__401__I
timestamp 1669390400
transform -1 0 26320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__402__I
timestamp 1669390400
transform 1 0 39984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A1
timestamp 1669390400
transform 1 0 42000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__403__A2
timestamp 1669390400
transform 1 0 41440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__405__I
timestamp 1669390400
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1669390400
transform -1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__408__I
timestamp 1669390400
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__409__I
timestamp 1669390400
transform 1 0 31024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A1
timestamp 1669390400
transform 1 0 34608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A2
timestamp 1669390400
transform -1 0 31024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__411__A3
timestamp 1669390400
transform 1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A1
timestamp 1669390400
transform 1 0 29680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__413__A2
timestamp 1669390400
transform -1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__414__I
timestamp 1669390400
transform 1 0 35840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__I
timestamp 1669390400
transform -1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A1
timestamp 1669390400
transform 1 0 35056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__419__A2
timestamp 1669390400
transform 1 0 35504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__420__I
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__I
timestamp 1669390400
transform 1 0 19488 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__I
timestamp 1669390400
transform -1 0 15568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A2
timestamp 1669390400
transform 1 0 15568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__I
timestamp 1669390400
transform 1 0 38528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A1
timestamp 1669390400
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A2
timestamp 1669390400
transform 1 0 36736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A3
timestamp 1669390400
transform 1 0 33488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__427__A4
timestamp 1669390400
transform -1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__429__I
timestamp 1669390400
transform 1 0 26992 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__430__B
timestamp 1669390400
transform 1 0 26544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A1
timestamp 1669390400
transform -1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__432__A2
timestamp 1669390400
transform 1 0 14448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A1
timestamp 1669390400
transform 1 0 15232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__433__A2
timestamp 1669390400
transform -1 0 15008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__434__A2
timestamp 1669390400
transform -1 0 5712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A2
timestamp 1669390400
transform -1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__437__B2
timestamp 1669390400
transform 1 0 7168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A2
timestamp 1669390400
transform 1 0 3472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__443__A2
timestamp 1669390400
transform 1 0 3136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__444__A1
timestamp 1669390400
transform 1 0 5264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__A2
timestamp 1669390400
transform 1 0 7616 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__B
timestamp 1669390400
transform 1 0 8064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__A2
timestamp 1669390400
transform 1 0 9184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__A2
timestamp 1669390400
transform -1 0 8736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__I
timestamp 1669390400
transform -1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__I
timestamp 1669390400
transform 1 0 27776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A1
timestamp 1669390400
transform 1 0 4368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__A2
timestamp 1669390400
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__A2
timestamp 1669390400
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__B
timestamp 1669390400
transform 1 0 11872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__A2
timestamp 1669390400
transform -1 0 11760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A1
timestamp 1669390400
transform 1 0 3584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__A2
timestamp 1669390400
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A1
timestamp 1669390400
transform -1 0 12544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__A2
timestamp 1669390400
transform 1 0 11984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__A1
timestamp 1669390400
transform 1 0 6048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A1
timestamp 1669390400
transform -1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A2
timestamp 1669390400
transform -1 0 11648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__A3
timestamp 1669390400
transform -1 0 2352 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__A1
timestamp 1669390400
transform 1 0 6384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__A2
timestamp 1669390400
transform 1 0 4480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__A2
timestamp 1669390400
transform -1 0 4256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A1
timestamp 1669390400
transform -1 0 3472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__A2
timestamp 1669390400
transform -1 0 1904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__B
timestamp 1669390400
transform -1 0 13104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A1
timestamp 1669390400
transform -1 0 11760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__A2
timestamp 1669390400
transform -1 0 11200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A1
timestamp 1669390400
transform 1 0 14224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__A2
timestamp 1669390400
transform 1 0 13328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__A2
timestamp 1669390400
transform 1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A1
timestamp 1669390400
transform -1 0 6384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__A2
timestamp 1669390400
transform 1 0 5712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__A2
timestamp 1669390400
transform -1 0 2800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__I
timestamp 1669390400
transform -1 0 12656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__A2
timestamp 1669390400
transform 1 0 15120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__A2
timestamp 1669390400
transform -1 0 1904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__B
timestamp 1669390400
transform -1 0 15456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A1
timestamp 1669390400
transform 1 0 4256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__A2
timestamp 1669390400
transform 1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A1
timestamp 1669390400
transform -1 0 3360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A2
timestamp 1669390400
transform -1 0 3808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__A3
timestamp 1669390400
transform -1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__A1
timestamp 1669390400
transform -1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__A2
timestamp 1669390400
transform 1 0 12880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__A1
timestamp 1669390400
transform -1 0 2352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A1
timestamp 1669390400
transform 1 0 18144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__A2
timestamp 1669390400
transform 1 0 19152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A1
timestamp 1669390400
transform -1 0 2576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__A2
timestamp 1669390400
transform -1 0 3136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__I
timestamp 1669390400
transform 1 0 9632 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__A1
timestamp 1669390400
transform -1 0 18368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__A2
timestamp 1669390400
transform -1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__A1
timestamp 1669390400
transform -1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A1
timestamp 1669390400
transform -1 0 16352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__A4
timestamp 1669390400
transform -1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__A2
timestamp 1669390400
transform -1 0 17696 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__A2
timestamp 1669390400
transform 1 0 2688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__A3
timestamp 1669390400
transform 1 0 16016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__A3
timestamp 1669390400
transform 1 0 17920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__A1
timestamp 1669390400
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__B
timestamp 1669390400
transform 1 0 32816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A1
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A2
timestamp 1669390400
transform 1 0 28672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A1
timestamp 1669390400
transform 1 0 25424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__A2
timestamp 1669390400
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__I
timestamp 1669390400
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__B2
timestamp 1669390400
transform -1 0 19264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A1
timestamp 1669390400
transform -1 0 2800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__503__A2
timestamp 1669390400
transform 1 0 17584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A1
timestamp 1669390400
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__A2
timestamp 1669390400
transform -1 0 17808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__B1
timestamp 1669390400
transform 1 0 28672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__504__C
timestamp 1669390400
transform -1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__A2
timestamp 1669390400
transform 1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__B1
timestamp 1669390400
transform -1 0 13888 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__B2
timestamp 1669390400
transform 1 0 38192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__505__C
timestamp 1669390400
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A1
timestamp 1669390400
transform -1 0 28112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__506__A2
timestamp 1669390400
transform -1 0 28560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A1
timestamp 1669390400
transform -1 0 27664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__507__A2
timestamp 1669390400
transform -1 0 27552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__508__A2
timestamp 1669390400
transform 1 0 33040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__510__A3
timestamp 1669390400
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A2
timestamp 1669390400
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__511__A3
timestamp 1669390400
transform 1 0 36512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__B1
timestamp 1669390400
transform -1 0 14112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__512__B2
timestamp 1669390400
transform 1 0 20832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A1
timestamp 1669390400
transform -1 0 34160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A2
timestamp 1669390400
transform -1 0 33488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1669390400
transform 1 0 16912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A2
timestamp 1669390400
transform 1 0 18704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A2
timestamp 1669390400
transform -1 0 18928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__515__A3
timestamp 1669390400
transform -1 0 26320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A1
timestamp 1669390400
transform 1 0 38416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__516__A2
timestamp 1669390400
transform 1 0 37408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A1
timestamp 1669390400
transform -1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A2
timestamp 1669390400
transform -1 0 16688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__517__A3
timestamp 1669390400
transform -1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__518__A2
timestamp 1669390400
transform -1 0 19936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A2
timestamp 1669390400
transform 1 0 42000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__B1
timestamp 1669390400
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__B2
timestamp 1669390400
transform 1 0 19936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__C
timestamp 1669390400
transform -1 0 7392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__B2
timestamp 1669390400
transform 1 0 19152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A1
timestamp 1669390400
transform 1 0 21280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__A2
timestamp 1669390400
transform 1 0 31248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__521__B
timestamp 1669390400
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A1
timestamp 1669390400
transform 1 0 37408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A2
timestamp 1669390400
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A1
timestamp 1669390400
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__523__A2
timestamp 1669390400
transform -1 0 22176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1669390400
transform -1 0 4144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A1
timestamp 1669390400
transform 1 0 20384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__525__A2
timestamp 1669390400
transform 1 0 20832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__526__A2
timestamp 1669390400
transform -1 0 29456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A1
timestamp 1669390400
transform -1 0 25872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__527__A2
timestamp 1669390400
transform -1 0 23072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A1
timestamp 1669390400
transform 1 0 34832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__528__A2
timestamp 1669390400
transform -1 0 32816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A2
timestamp 1669390400
transform 1 0 29232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__A3
timestamp 1669390400
transform 1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__A2
timestamp 1669390400
transform 1 0 25536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__B1
timestamp 1669390400
transform 1 0 26432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__B2
timestamp 1669390400
transform 1 0 24640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__530__C
timestamp 1669390400
transform -1 0 27664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__531__I
timestamp 1669390400
transform -1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__B1
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__532__B2
timestamp 1669390400
transform 1 0 24192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A1
timestamp 1669390400
transform -1 0 38416 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__533__A2
timestamp 1669390400
transform -1 0 38864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__534__I
timestamp 1669390400
transform 1 0 30800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__A1
timestamp 1669390400
transform 1 0 33936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__A2
timestamp 1669390400
transform 1 0 39648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A1
timestamp 1669390400
transform -1 0 30128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__A2
timestamp 1669390400
transform 1 0 31696 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__537__B
timestamp 1669390400
transform -1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A1
timestamp 1669390400
transform 1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__538__A2
timestamp 1669390400
transform -1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__A2
timestamp 1669390400
transform -1 0 18816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B1
timestamp 1669390400
transform -1 0 27216 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__B2
timestamp 1669390400
transform -1 0 3248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__539__C
timestamp 1669390400
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B1
timestamp 1669390400
transform -1 0 21728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__540__B2
timestamp 1669390400
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__A1
timestamp 1669390400
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__541__B
timestamp 1669390400
transform -1 0 26320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__543__A1
timestamp 1669390400
transform 1 0 28784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A1
timestamp 1669390400
transform 1 0 31248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__544__A2
timestamp 1669390400
transform 1 0 31360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__545__I
timestamp 1669390400
transform 1 0 32144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A1
timestamp 1669390400
transform 1 0 33712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__546__A2
timestamp 1669390400
transform -1 0 31248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A1
timestamp 1669390400
transform -1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__548__A2
timestamp 1669390400
transform -1 0 31024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A1
timestamp 1669390400
transform 1 0 39872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__549__A2
timestamp 1669390400
transform 1 0 35728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__A2
timestamp 1669390400
transform 1 0 32144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__550__A3
timestamp 1669390400
transform -1 0 31472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__A2
timestamp 1669390400
transform -1 0 30240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__B1
timestamp 1669390400
transform -1 0 31920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__B2
timestamp 1669390400
transform -1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__551__C
timestamp 1669390400
transform -1 0 33040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__552__I
timestamp 1669390400
transform 1 0 35056 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__B1
timestamp 1669390400
transform 1 0 38304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__553__B2
timestamp 1669390400
transform -1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__A1
timestamp 1669390400
transform 1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__554__A2
timestamp 1669390400
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A1
timestamp 1669390400
transform 1 0 37856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__555__A2
timestamp 1669390400
transform 1 0 38864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__556__I
timestamp 1669390400
transform 1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A1
timestamp 1669390400
transform 1 0 35952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__557__A2
timestamp 1669390400
transform -1 0 36848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A1
timestamp 1669390400
transform -1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__558__A2
timestamp 1669390400
transform 1 0 32592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A1
timestamp 1669390400
transform 1 0 37856 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__559__A2
timestamp 1669390400
transform 1 0 38864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A1
timestamp 1669390400
transform -1 0 32592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A2
timestamp 1669390400
transform -1 0 31696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__560__A3
timestamp 1669390400
transform -1 0 33040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__561__A2
timestamp 1669390400
transform 1 0 31920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__A2
timestamp 1669390400
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B1
timestamp 1669390400
transform -1 0 34832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B2
timestamp 1669390400
transform 1 0 38976 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__C
timestamp 1669390400
transform -1 0 32144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__563__I
timestamp 1669390400
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B1
timestamp 1669390400
transform -1 0 32592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__B2
timestamp 1669390400
transform 1 0 39424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A1
timestamp 1669390400
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__565__A2
timestamp 1669390400
transform 1 0 37520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A1
timestamp 1669390400
transform 1 0 39200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__566__A2
timestamp 1669390400
transform 1 0 38416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A1
timestamp 1669390400
transform -1 0 30576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__567__A2
timestamp 1669390400
transform -1 0 30576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1669390400
transform -1 0 28000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__569__I
timestamp 1669390400
transform 1 0 40992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A1
timestamp 1669390400
transform 1 0 33600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__570__A2
timestamp 1669390400
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__571__B
timestamp 1669390400
transform -1 0 31136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__A1
timestamp 1669390400
transform -1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__572__A2
timestamp 1669390400
transform -1 0 41888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__A1
timestamp 1669390400
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__574__A2
timestamp 1669390400
transform 1 0 41216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A1
timestamp 1669390400
transform 1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__575__A2
timestamp 1669390400
transform 1 0 40208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__578__I
timestamp 1669390400
transform -1 0 41776 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A1
timestamp 1669390400
transform -1 0 38752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__580__A2
timestamp 1669390400
transform -1 0 38304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__A2
timestamp 1669390400
transform 1 0 39312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__B1
timestamp 1669390400
transform 1 0 39312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__B2
timestamp 1669390400
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__581__C
timestamp 1669390400
transform 1 0 39760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__B1
timestamp 1669390400
transform -1 0 39200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__582__B2
timestamp 1669390400
transform -1 0 36960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__583__A1
timestamp 1669390400
transform 1 0 42000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A1
timestamp 1669390400
transform 1 0 41888 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__A2
timestamp 1669390400
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__585__A1
timestamp 1669390400
transform -1 0 41776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__586__I
timestamp 1669390400
transform 1 0 42000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A1
timestamp 1669390400
transform -1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__A2
timestamp 1669390400
transform -1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__587__B
timestamp 1669390400
transform 1 0 20832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A1
timestamp 1669390400
transform -1 0 23072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__588__A2
timestamp 1669390400
transform -1 0 18704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__A2
timestamp 1669390400
transform -1 0 35952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__B1
timestamp 1669390400
transform -1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__589__C
timestamp 1669390400
transform 1 0 36176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__B1
timestamp 1669390400
transform -1 0 37744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__B2
timestamp 1669390400
transform -1 0 35840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__591__A2
timestamp 1669390400
transform -1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__A2
timestamp 1669390400
transform 1 0 42000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A2
timestamp 1669390400
transform 1 0 42000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A2
timestamp 1669390400
transform -1 0 37856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A1
timestamp 1669390400
transform 1 0 37408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A2
timestamp 1669390400
transform -1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__B1
timestamp 1669390400
transform -1 0 35504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__C
timestamp 1669390400
transform 1 0 34832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__601__B2
timestamp 1669390400
transform 1 0 37520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1669390400
transform -1 0 41440 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__603__A1
timestamp 1669390400
transform 1 0 40992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A2
timestamp 1669390400
transform 1 0 39984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A1
timestamp 1669390400
transform -1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A2
timestamp 1669390400
transform 1 0 37856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__B1
timestamp 1669390400
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__C
timestamp 1669390400
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__B1
timestamp 1669390400
transform 1 0 37408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__609__B2
timestamp 1669390400
transform -1 0 33712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A1
timestamp 1669390400
transform 1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__612__A2
timestamp 1669390400
transform 1 0 40432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__617__A2
timestamp 1669390400
transform 1 0 38304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A1
timestamp 1669390400
transform 1 0 40432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__618__A2
timestamp 1669390400
transform 1 0 39984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__622__A2
timestamp 1669390400
transform 1 0 39200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__A2
timestamp 1669390400
transform 1 0 34832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__B1
timestamp 1669390400
transform 1 0 35728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__B2
timestamp 1669390400
transform 1 0 37968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__623__C
timestamp 1669390400
transform 1 0 35280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__624__B2
timestamp 1669390400
transform 1 0 33936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__627__A2
timestamp 1669390400
transform 1 0 36176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__628__A1
timestamp 1669390400
transform 1 0 37072 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__A3
timestamp 1669390400
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__A2
timestamp 1669390400
transform 1 0 34384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__B1
timestamp 1669390400
transform 1 0 34384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__B2
timestamp 1669390400
transform -1 0 35504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__632__C
timestamp 1669390400
transform 1 0 35728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__633__B2
timestamp 1669390400
transform 1 0 37744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__645__A2
timestamp 1669390400
transform 1 0 38080 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A1
timestamp 1669390400
transform -1 0 35504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__A2
timestamp 1669390400
transform 1 0 33488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__B1
timestamp 1669390400
transform 1 0 33936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__B2
timestamp 1669390400
transform -1 0 36848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__C
timestamp 1669390400
transform 1 0 34384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__647__B2
timestamp 1669390400
transform 1 0 32256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__650__A1
timestamp 1669390400
transform 1 0 34160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__651__A1
timestamp 1669390400
transform 1 0 36176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__655__A3
timestamp 1669390400
transform 1 0 35728 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A1
timestamp 1669390400
transform -1 0 30576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__A2
timestamp 1669390400
transform 1 0 28672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__B1
timestamp 1669390400
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__B2
timestamp 1669390400
transform -1 0 31920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__656__C
timestamp 1669390400
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A1
timestamp 1669390400
transform 1 0 38080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__657__A2
timestamp 1669390400
transform -1 0 30240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__658__A1
timestamp 1669390400
transform 1 0 39984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__A1
timestamp 1669390400
transform -1 0 34160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__A2
timestamp 1669390400
transform -1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__A1
timestamp 1669390400
transform 1 0 30464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__A2
timestamp 1669390400
transform -1 0 31136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A1
timestamp 1669390400
transform -1 0 33040 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__A2
timestamp 1669390400
transform -1 0 32928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A1
timestamp 1669390400
transform 1 0 27776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__A2
timestamp 1669390400
transform 1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A1
timestamp 1669390400
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__A2
timestamp 1669390400
transform 1 0 31808 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__B1
timestamp 1669390400
transform -1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__B2
timestamp 1669390400
transform 1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__B
timestamp 1669390400
transform 1 0 28112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__A1
timestamp 1669390400
transform 1 0 31920 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__A2
timestamp 1669390400
transform 1 0 31584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A1
timestamp 1669390400
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__A2
timestamp 1669390400
transform -1 0 28000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__B2
timestamp 1669390400
transform 1 0 21728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__687__B
timestamp 1669390400
transform -1 0 26656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A1
timestamp 1669390400
transform 1 0 29904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__A2
timestamp 1669390400
transform 1 0 31472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__B
timestamp 1669390400
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__691__A2
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__692__A2
timestamp 1669390400
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__A1
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__B2
timestamp 1669390400
transform 1 0 22960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__699__B
timestamp 1669390400
transform 1 0 22176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A1
timestamp 1669390400
transform 1 0 26320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__705__A1
timestamp 1669390400
transform 1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__707__CLK
timestamp 1669390400
transform -1 0 14000 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__CLK
timestamp 1669390400
transform 1 0 10080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__709__CLK
timestamp 1669390400
transform 1 0 1904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__710__CLK
timestamp 1669390400
transform -1 0 5152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__CLK
timestamp 1669390400
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__712__CLK
timestamp 1669390400
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__713__CLK
timestamp 1669390400
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__714__CLK
timestamp 1669390400
transform 1 0 4144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__715__CLK
timestamp 1669390400
transform 1 0 3024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__CLK
timestamp 1669390400
transform -1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__717__CLK
timestamp 1669390400
transform 1 0 4704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__718__CLK
timestamp 1669390400
transform -1 0 2016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__719__CLK
timestamp 1669390400
transform 1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__720__CLK
timestamp 1669390400
transform 1 0 16464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__721__CLK
timestamp 1669390400
transform 1 0 14672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__722__CLK
timestamp 1669390400
transform -1 0 15904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__CLK
timestamp 1669390400
transform 1 0 35392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__724__CLK
timestamp 1669390400
transform -1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__725__CLK
timestamp 1669390400
transform -1 0 16464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__726__CLK
timestamp 1669390400
transform 1 0 18256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__727__CLK
timestamp 1669390400
transform 1 0 23296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__728__CLK
timestamp 1669390400
transform 1 0 26544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__729__CLK
timestamp 1669390400
transform 1 0 25536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__CLK
timestamp 1669390400
transform 1 0 33488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__CLK
timestamp 1669390400
transform -1 0 33936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__CLK
timestamp 1669390400
transform 1 0 37072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__CLK
timestamp 1669390400
transform 1 0 34160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__734__CLK
timestamp 1669390400
transform 1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__735__CLK
timestamp 1669390400
transform -1 0 32368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__CLK
timestamp 1669390400
transform 1 0 33488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__737__CLK
timestamp 1669390400
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__CLK
timestamp 1669390400
transform 1 0 28672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__CLK
timestamp 1669390400
transform 1 0 26656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__CLK
timestamp 1669390400
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__741__CLK
timestamp 1669390400
transform 1 0 25872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__CLK
timestamp 1669390400
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__743__CLK
timestamp 1669390400
transform 1 0 20832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__744__CLK
timestamp 1669390400
transform 1 0 16912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1669390400
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1669390400
transform 1 0 16912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1669390400
transform -1 0 28672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1669390400
transform 1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 3696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 39424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 22176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 35392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 40320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 40768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 19600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform -1 0 24416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform -1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform -1 0 23968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 33264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform 1 0 40544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform 1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform -1 0 20160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform -1 0 1904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 38304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1669390400
transform -1 0 15344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1669390400
transform -1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18
timestamp 1669390400
transform 1 0 3360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53
timestamp 1669390400
transform 1 0 7280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1669390400
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122
timestamp 1669390400
transform 1 0 15008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_124
timestamp 1669390400
transform 1 0 15232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_158
timestamp 1669390400
transform 1 0 19040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_182
timestamp 1669390400
transform 1 0 21728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_229
timestamp 1669390400
transform 1 0 26992 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1669390400
transform 1 0 28224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_264 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30912 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_299
timestamp 1669390400
transform 1 0 34832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_311
timestamp 1669390400
transform 1 0 36176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_334
timestamp 1669390400
transform 1 0 38752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_344
timestamp 1669390400
transform 1 0 39872 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_348
timestamp 1669390400
transform 1 0 40320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_361
timestamp 1669390400
transform 1 0 41776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_365
timestamp 1669390400
transform 1 0 42224 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_17
timestamp 1669390400
transform 1 0 3248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_25
timestamp 1669390400
transform 1 0 4144 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_33
timestamp 1669390400
transform 1 0 5040 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_49
timestamp 1669390400
transform 1 0 6832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_51
timestamp 1669390400
transform 1 0 7056 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1669390400
transform 1 0 7392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_103
timestamp 1669390400
transform 1 0 12880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_107
timestamp 1669390400
transform 1 0 13328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_117
timestamp 1669390400
transform 1 0 14448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_133
timestamp 1669390400
transform 1 0 16240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_175
timestamp 1669390400
transform 1 0 20944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_206
timestamp 1669390400
transform 1 0 24416 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_221
timestamp 1669390400
transform 1 0 26096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_252
timestamp 1669390400
transform 1 0 29568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_316
timestamp 1669390400
transform 1 0 36736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_334
timestamp 1669390400
transform 1 0 38752 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_352
timestamp 1669390400
transform 1 0 40768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_364
timestamp 1669390400
transform 1 0 42112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_8
timestamp 1669390400
transform 1 0 2240 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_12
timestamp 1669390400
transform 1 0 2688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_18
timestamp 1669390400
transform 1 0 3360 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_20
timestamp 1669390400
transform 1 0 3584 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_26
timestamp 1669390400
transform 1 0 4256 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_46
timestamp 1669390400
transform 1 0 6496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_77
timestamp 1669390400
transform 1 0 9968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_81
timestamp 1669390400
transform 1 0 10416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_91
timestamp 1669390400
transform 1 0 11536 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_112
timestamp 1669390400
transform 1 0 13888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_143
timestamp 1669390400
transform 1 0 17360 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_159
timestamp 1669390400
transform 1 0 19152 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_166
timestamp 1669390400
transform 1 0 19936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_194
timestamp 1669390400
transform 1 0 23072 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_196
timestamp 1669390400
transform 1 0 23296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_207
timestamp 1669390400
transform 1 0 24528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_213
timestamp 1669390400
transform 1 0 25200 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_231
timestamp 1669390400
transform 1 0 27216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_235
timestamp 1669390400
transform 1 0 27664 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_267
timestamp 1669390400
transform 1 0 31248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_285
timestamp 1669390400
transform 1 0 33264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_303
timestamp 1669390400
transform 1 0 35280 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_315
timestamp 1669390400
transform 1 0 36624 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_339
timestamp 1669390400
transform 1 0 39312 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_357
timestamp 1669390400
transform 1 0 41328 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_5
timestamp 1669390400
transform 1 0 1904 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_9
timestamp 1669390400
transform 1 0 2352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_13
timestamp 1669390400
transform 1 0 2800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_17
timestamp 1669390400
transform 1 0 3248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_21
timestamp 1669390400
transform 1 0 3696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_25
timestamp 1669390400
transform 1 0 4144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_33
timestamp 1669390400
transform 1 0 5040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_41
timestamp 1669390400
transform 1 0 5936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_52
timestamp 1669390400
transform 1 0 7168 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_64
timestamp 1669390400
transform 1 0 8512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1669390400
transform 1 0 9856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_84
timestamp 1669390400
transform 1 0 10752 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_94
timestamp 1669390400
transform 1 0 11872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_109
timestamp 1669390400
transform 1 0 13552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_111
timestamp 1669390400
transform 1 0 13776 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_114
timestamp 1669390400
transform 1 0 14112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_124
timestamp 1669390400
transform 1 0 15232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_134
timestamp 1669390400
transform 1 0 16352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_162
timestamp 1669390400
transform 1 0 19488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_166
timestamp 1669390400
transform 1 0 19936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_197
timestamp 1669390400
transform 1 0 23408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_218
timestamp 1669390400
transform 1 0 25760 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_231
timestamp 1669390400
transform 1 0 27216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_237
timestamp 1669390400
transform 1 0 27888 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_255
timestamp 1669390400
transform 1 0 29904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_259
timestamp 1669390400
transform 1 0 30352 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_271
timestamp 1669390400
transform 1 0 31696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_316
timestamp 1669390400
transform 1 0 36736 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_327
timestamp 1669390400
transform 1 0 37968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_331
timestamp 1669390400
transform 1 0 38416 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_333
timestamp 1669390400
transform 1 0 38640 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_363
timestamp 1669390400
transform 1 0 42000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_365
timestamp 1669390400
transform 1 0 42224 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1669390400
transform 1 0 2016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_10
timestamp 1669390400
transform 1 0 2464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1669390400
transform 1 0 2912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_18
timestamp 1669390400
transform 1 0 3360 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_22
timestamp 1669390400
transform 1 0 3808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_28
timestamp 1669390400
transform 1 0 4480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_43
timestamp 1669390400
transform 1 0 6160 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_74
timestamp 1669390400
transform 1 0 9632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_110
timestamp 1669390400
transform 1 0 13664 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_140
timestamp 1669390400
transform 1 0 17024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_149
timestamp 1669390400
transform 1 0 18032 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_159
timestamp 1669390400
transform 1 0 19152 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_169
timestamp 1669390400
transform 1 0 20272 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_188
timestamp 1669390400
transform 1 0 22400 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_199
timestamp 1669390400
transform 1 0 23632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_210
timestamp 1669390400
transform 1 0 24864 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_221
timestamp 1669390400
transform 1 0 26096 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_231
timestamp 1669390400
transform 1 0 27216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_241
timestamp 1669390400
transform 1 0 28336 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_261
timestamp 1669390400
transform 1 0 30576 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_272
timestamp 1669390400
transform 1 0 31808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_303
timestamp 1669390400
transform 1 0 35280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_307
timestamp 1669390400
transform 1 0 35728 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_317
timestamp 1669390400
transform 1 0 36848 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_332
timestamp 1669390400
transform 1 0 38528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_350
timestamp 1669390400
transform 1 0 40544 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_357
timestamp 1669390400
transform 1 0 41328 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_364
timestamp 1669390400
transform 1 0 42112 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_5
timestamp 1669390400
transform 1 0 1904 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_9
timestamp 1669390400
transform 1 0 2352 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_13
timestamp 1669390400
transform 1 0 2800 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_17
timestamp 1669390400
transform 1 0 3248 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_23
timestamp 1669390400
transform 1 0 3920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_29
timestamp 1669390400
transform 1 0 4592 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_36
timestamp 1669390400
transform 1 0 5376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_43
timestamp 1669390400
transform 1 0 6160 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_54
timestamp 1669390400
transform 1 0 7392 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_60
timestamp 1669390400
transform 1 0 8064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_86
timestamp 1669390400
transform 1 0 10976 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_140
timestamp 1669390400
transform 1 0 17024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_174
timestamp 1669390400
transform 1 0 20832 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_182
timestamp 1669390400
transform 1 0 21728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_190
timestamp 1669390400
transform 1 0 22624 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_203
timestamp 1669390400
transform 1 0 24080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1669390400
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_218
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_220
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_229
timestamp 1669390400
transform 1 0 26992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_239
timestamp 1669390400
transform 1 0 28112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_249
timestamp 1669390400
transform 1 0 29232 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_257
timestamp 1669390400
transform 1 0 30128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_265
timestamp 1669390400
transform 1 0 31024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_269
timestamp 1669390400
transform 1 0 31472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1669390400
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_293
timestamp 1669390400
transform 1 0 34160 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_295
timestamp 1669390400
transform 1 0 34384 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_307
timestamp 1669390400
transform 1 0 35728 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_320
timestamp 1669390400
transform 1 0 37184 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_324
timestamp 1669390400
transform 1 0 37632 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_333
timestamp 1669390400
transform 1 0 38640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_341
timestamp 1669390400
transform 1 0 39536 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_349
timestamp 1669390400
transform 1 0 40432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_353
timestamp 1669390400
transform 1 0 40880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_363
timestamp 1669390400
transform 1 0 42000 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_365
timestamp 1669390400
transform 1 0 42224 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_4
timestamp 1669390400
transform 1 0 1792 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_7
timestamp 1669390400
transform 1 0 2128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_11
timestamp 1669390400
transform 1 0 2576 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_15
timestamp 1669390400
transform 1 0 3024 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_19
timestamp 1669390400
transform 1 0 3472 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_23
timestamp 1669390400
transform 1 0 3920 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_27
timestamp 1669390400
transform 1 0 4368 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_43
timestamp 1669390400
transform 1 0 6160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_51
timestamp 1669390400
transform 1 0 7056 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_58
timestamp 1669390400
transform 1 0 7840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_66
timestamp 1669390400
transform 1 0 8736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_74
timestamp 1669390400
transform 1 0 9632 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_116
timestamp 1669390400
transform 1 0 14336 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_126
timestamp 1669390400
transform 1 0 15456 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_159
timestamp 1669390400
transform 1 0 19152 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_161
timestamp 1669390400
transform 1 0 19376 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_168
timestamp 1669390400
transform 1 0 20160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_190
timestamp 1669390400
transform 1 0 22624 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1669390400
transform 1 0 28448 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_246
timestamp 1669390400
transform 1 0 28896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_257
timestamp 1669390400
transform 1 0 30128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_265
timestamp 1669390400
transform 1 0 31024 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_273
timestamp 1669390400
transform 1 0 31920 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_277
timestamp 1669390400
transform 1 0 32368 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_307
timestamp 1669390400
transform 1 0 35728 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_327
timestamp 1669390400
transform 1 0 37968 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_329
timestamp 1669390400
transform 1 0 38192 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_338
timestamp 1669390400
transform 1 0 39200 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_348
timestamp 1669390400
transform 1 0 40320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_356
timestamp 1669390400
transform 1 0 41216 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_363
timestamp 1669390400
transform 1 0 42000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_365
timestamp 1669390400
transform 1 0 42224 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_8
timestamp 1669390400
transform 1 0 2240 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_12
timestamp 1669390400
transform 1 0 2688 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_16
timestamp 1669390400
transform 1 0 3136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_20
timestamp 1669390400
transform 1 0 3584 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_24
timestamp 1669390400
transform 1 0 4032 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_28
timestamp 1669390400
transform 1 0 4480 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_32
timestamp 1669390400
transform 1 0 4928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1669390400
transform 1 0 5600 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_45
timestamp 1669390400
transform 1 0 6384 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_52
timestamp 1669390400
transform 1 0 7168 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_62
timestamp 1669390400
transform 1 0 8288 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_80
timestamp 1669390400
transform 1 0 10304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_88
timestamp 1669390400
transform 1 0 11200 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_140
timestamp 1669390400
transform 1 0 17024 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_147
timestamp 1669390400
transform 1 0 17808 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_155
timestamp 1669390400
transform 1 0 18704 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_157
timestamp 1669390400
transform 1 0 18928 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1669390400
transform 1 0 19264 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_191
timestamp 1669390400
transform 1 0 22736 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_201
timestamp 1669390400
transform 1 0 23856 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_211
timestamp 1669390400
transform 1 0 24976 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_223
timestamp 1669390400
transform 1 0 26320 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_232
timestamp 1669390400
transform 1 0 27328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_239
timestamp 1669390400
transform 1 0 28112 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_249
timestamp 1669390400
transform 1 0 29232 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_257
timestamp 1669390400
transform 1 0 30128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_261
timestamp 1669390400
transform 1 0 30576 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_269
timestamp 1669390400
transform 1 0 31472 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_278
timestamp 1669390400
transform 1 0 32480 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_282
timestamp 1669390400
transform 1 0 32928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_293
timestamp 1669390400
transform 1 0 34160 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_301
timestamp 1669390400
transform 1 0 35056 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_309
timestamp 1669390400
transform 1 0 35952 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_317
timestamp 1669390400
transform 1 0 36848 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_324
timestamp 1669390400
transform 1 0 37632 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_331
timestamp 1669390400
transform 1 0 38416 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_338
timestamp 1669390400
transform 1 0 39200 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_345
timestamp 1669390400
transform 1 0 39984 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_352
timestamp 1669390400
transform 1 0 40768 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_363
timestamp 1669390400
transform 1 0 42000 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_365
timestamp 1669390400
transform 1 0 42224 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1669390400
transform 1 0 2016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_10
timestamp 1669390400
transform 1 0 2464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_14
timestamp 1669390400
transform 1 0 2912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_18
timestamp 1669390400
transform 1 0 3360 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_22
timestamp 1669390400
transform 1 0 3808 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_26
timestamp 1669390400
transform 1 0 4256 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_30
timestamp 1669390400
transform 1 0 4704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_40
timestamp 1669390400
transform 1 0 5824 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_44
timestamp 1669390400
transform 1 0 6272 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_75
timestamp 1669390400
transform 1 0 9744 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_83
timestamp 1669390400
transform 1 0 10640 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_95
timestamp 1669390400
transform 1 0 11984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_138
timestamp 1669390400
transform 1 0 16800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_148
timestamp 1669390400
transform 1 0 17920 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_155
timestamp 1669390400
transform 1 0 18704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_165
timestamp 1669390400
transform 1 0 19824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_169
timestamp 1669390400
transform 1 0 20272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_192
timestamp 1669390400
transform 1 0 22848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_196
timestamp 1669390400
transform 1 0 23296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_204
timestamp 1669390400
transform 1 0 24192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_213
timestamp 1669390400
transform 1 0 25200 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_217
timestamp 1669390400
transform 1 0 25648 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_219
timestamp 1669390400
transform 1 0 25872 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_228
timestamp 1669390400
transform 1 0 26880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_238
timestamp 1669390400
transform 1 0 28000 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_253
timestamp 1669390400
transform 1 0 29680 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_263
timestamp 1669390400
transform 1 0 30800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_272
timestamp 1669390400
transform 1 0 31808 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_305
timestamp 1669390400
transform 1 0 35504 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_312
timestamp 1669390400
transform 1 0 36288 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_329
timestamp 1669390400
transform 1 0 38192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_337
timestamp 1669390400
transform 1 0 39088 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_339
timestamp 1669390400
transform 1 0 39312 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_348
timestamp 1669390400
transform 1 0 40320 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_355
timestamp 1669390400
transform 1 0 41104 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_362
timestamp 1669390400
transform 1 0 41888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_10
timestamp 1669390400
transform 1 0 2464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_13
timestamp 1669390400
transform 1 0 2800 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_17
timestamp 1669390400
transform 1 0 3248 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_21
timestamp 1669390400
transform 1 0 3696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_25
timestamp 1669390400
transform 1 0 4144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_29
timestamp 1669390400
transform 1 0 4592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_33
timestamp 1669390400
transform 1 0 5040 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_37
timestamp 1669390400
transform 1 0 5488 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_41
timestamp 1669390400
transform 1 0 5936 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_45
timestamp 1669390400
transform 1 0 6384 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_51
timestamp 1669390400
transform 1 0 7056 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_59
timestamp 1669390400
transform 1 0 7952 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_79
timestamp 1669390400
transform 1 0 10192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_83
timestamp 1669390400
transform 1 0 10640 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_113
timestamp 1669390400
transform 1 0 14000 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_121
timestamp 1669390400
transform 1 0 14896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_131
timestamp 1669390400
transform 1 0 16016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_152
timestamp 1669390400
transform 1 0 18368 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_160
timestamp 1669390400
transform 1 0 19264 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_164
timestamp 1669390400
transform 1 0 19712 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_194
timestamp 1669390400
transform 1 0 23072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_200
timestamp 1669390400
transform 1 0 23744 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_211
timestamp 1669390400
transform 1 0 24976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_229
timestamp 1669390400
transform 1 0 26992 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_239
timestamp 1669390400
transform 1 0 28112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_246
timestamp 1669390400
transform 1 0 28896 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_256
timestamp 1669390400
transform 1 0 30016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_264
timestamp 1669390400
transform 1 0 30912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_271
timestamp 1669390400
transform 1 0 31696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1669390400
transform 1 0 32928 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_292
timestamp 1669390400
transform 1 0 34048 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_305
timestamp 1669390400
transform 1 0 35504 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_312
timestamp 1669390400
transform 1 0 36288 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_316
timestamp 1669390400
transform 1 0 36736 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_326
timestamp 1669390400
transform 1 0 37856 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_336
timestamp 1669390400
transform 1 0 38976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_345
timestamp 1669390400
transform 1 0 39984 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_363
timestamp 1669390400
transform 1 0 42000 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_365
timestamp 1669390400
transform 1 0 42224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_18
timestamp 1669390400
transform 1 0 3360 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_22
timestamp 1669390400
transform 1 0 3808 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_26
timestamp 1669390400
transform 1 0 4256 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_30
timestamp 1669390400
transform 1 0 4704 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_45
timestamp 1669390400
transform 1 0 6384 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1669390400
transform 1 0 7280 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_63
timestamp 1669390400
transform 1 0 8400 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_70
timestamp 1669390400
transform 1 0 9184 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_72
timestamp 1669390400
transform 1 0 9408 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_79
timestamp 1669390400
transform 1 0 10192 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_83
timestamp 1669390400
transform 1 0 10640 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_89
timestamp 1669390400
transform 1 0 11312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_99
timestamp 1669390400
transform 1 0 12432 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_116
timestamp 1669390400
transform 1 0 14336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_122
timestamp 1669390400
transform 1 0 15008 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_132
timestamp 1669390400
transform 1 0 16128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_163
timestamp 1669390400
transform 1 0 19600 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_173
timestamp 1669390400
transform 1 0 20720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_190
timestamp 1669390400
transform 1 0 22624 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_242
timestamp 1669390400
transform 1 0 28448 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_246
timestamp 1669390400
transform 1 0 28896 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_260
timestamp 1669390400
transform 1 0 30464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_270
timestamp 1669390400
transform 1 0 31584 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_278
timestamp 1669390400
transform 1 0 32480 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_285
timestamp 1669390400
transform 1 0 33264 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_289
timestamp 1669390400
transform 1 0 33712 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_291
timestamp 1669390400
transform 1 0 33936 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_303
timestamp 1669390400
transform 1 0 35280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_307
timestamp 1669390400
transform 1 0 35728 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_327
timestamp 1669390400
transform 1 0 37968 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_334
timestamp 1669390400
transform 1 0 38752 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_338
timestamp 1669390400
transform 1 0 39200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_345
timestamp 1669390400
transform 1 0 39984 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_352
timestamp 1669390400
transform 1 0 40768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_359
timestamp 1669390400
transform 1 0 41552 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_365
timestamp 1669390400
transform 1 0 42224 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_18
timestamp 1669390400
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_26
timestamp 1669390400
transform 1 0 4256 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_28
timestamp 1669390400
transform 1 0 4480 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_31
timestamp 1669390400
transform 1 0 4816 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_35
timestamp 1669390400
transform 1 0 5264 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_39
timestamp 1669390400
transform 1 0 5712 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_83
timestamp 1669390400
transform 1 0 10640 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_89
timestamp 1669390400
transform 1 0 11312 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_91
timestamp 1669390400
transform 1 0 11536 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_98
timestamp 1669390400
transform 1 0 12320 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_105
timestamp 1669390400
transform 1 0 13104 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_112
timestamp 1669390400
transform 1 0 13888 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_119
timestamp 1669390400
transform 1 0 14672 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_126
timestamp 1669390400
transform 1 0 15456 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_128
timestamp 1669390400
transform 1 0 15680 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_131
timestamp 1669390400
transform 1 0 16016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_135
timestamp 1669390400
transform 1 0 16464 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_147
timestamp 1669390400
transform 1 0 17808 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_153
timestamp 1669390400
transform 1 0 18480 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_160
timestamp 1669390400
transform 1 0 19264 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_221
timestamp 1669390400
transform 1 0 26096 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_223
timestamp 1669390400
transform 1 0 26320 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_236
timestamp 1669390400
transform 1 0 27776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_243
timestamp 1669390400
transform 1 0 28560 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_256
timestamp 1669390400
transform 1 0 30016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_258
timestamp 1669390400
transform 1 0 30240 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_269
timestamp 1669390400
transform 1 0 31472 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_298
timestamp 1669390400
transform 1 0 34720 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_311
timestamp 1669390400
transform 1 0 36176 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_318
timestamp 1669390400
transform 1 0 36960 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_325
timestamp 1669390400
transform 1 0 37744 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_327
timestamp 1669390400
transform 1 0 37968 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_335
timestamp 1669390400
transform 1 0 38864 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_345
timestamp 1669390400
transform 1 0 39984 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_352
timestamp 1669390400
transform 1 0 40768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_363
timestamp 1669390400
transform 1 0 42000 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_365
timestamp 1669390400
transform 1 0 42224 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_43
timestamp 1669390400
transform 1 0 6160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_47
timestamp 1669390400
transform 1 0 6608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_80
timestamp 1669390400
transform 1 0 10304 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_86
timestamp 1669390400
transform 1 0 10976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_92
timestamp 1669390400
transform 1 0 11648 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_98
timestamp 1669390400
transform 1 0 12320 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_104
timestamp 1669390400
transform 1 0 12992 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_114
timestamp 1669390400
transform 1 0 14112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_120
timestamp 1669390400
transform 1 0 14784 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_124
timestamp 1669390400
transform 1 0 15232 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_127
timestamp 1669390400
transform 1 0 15568 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_131
timestamp 1669390400
transform 1 0 16016 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_135
timestamp 1669390400
transform 1 0 16464 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_139
timestamp 1669390400
transform 1 0 16912 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_143
timestamp 1669390400
transform 1 0 17360 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_149
timestamp 1669390400
transform 1 0 18032 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_155
timestamp 1669390400
transform 1 0 18704 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_159
timestamp 1669390400
transform 1 0 19152 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_166
timestamp 1669390400
transform 1 0 19936 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_189
timestamp 1669390400
transform 1 0 22512 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_199
timestamp 1669390400
transform 1 0 23632 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_232
timestamp 1669390400
transform 1 0 27328 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_259
timestamp 1669390400
transform 1 0 30352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_266
timestamp 1669390400
transform 1 0 31136 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_273
timestamp 1669390400
transform 1 0 31920 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_304
timestamp 1669390400
transform 1 0 35392 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_311
timestamp 1669390400
transform 1 0 36176 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_331
timestamp 1669390400
transform 1 0 38416 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_340
timestamp 1669390400
transform 1 0 39424 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_347
timestamp 1669390400
transform 1 0 40208 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_354
timestamp 1669390400
transform 1 0 40992 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_363
timestamp 1669390400
transform 1 0 42000 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_365
timestamp 1669390400
transform 1 0 42224 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_34
timestamp 1669390400
transform 1 0 5152 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_42
timestamp 1669390400
transform 1 0 6048 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_46
timestamp 1669390400
transform 1 0 6496 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_50
timestamp 1669390400
transform 1 0 6944 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_54
timestamp 1669390400
transform 1 0 7392 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_58
timestamp 1669390400
transform 1 0 7840 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_62
timestamp 1669390400
transform 1 0 8288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_75
timestamp 1669390400
transform 1 0 9744 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_78
timestamp 1669390400
transform 1 0 10080 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_82
timestamp 1669390400
transform 1 0 10528 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_86
timestamp 1669390400
transform 1 0 10976 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_89
timestamp 1669390400
transform 1 0 11312 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_93
timestamp 1669390400
transform 1 0 11760 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_97
timestamp 1669390400
transform 1 0 12208 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_101
timestamp 1669390400
transform 1 0 12656 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_105
timestamp 1669390400
transform 1 0 13104 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_109
timestamp 1669390400
transform 1 0 13552 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_113
timestamp 1669390400
transform 1 0 14000 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_117
timestamp 1669390400
transform 1 0 14448 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_121
timestamp 1669390400
transform 1 0 14896 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_125
timestamp 1669390400
transform 1 0 15344 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_129
timestamp 1669390400
transform 1 0 15792 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_133
timestamp 1669390400
transform 1 0 16240 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_175
timestamp 1669390400
transform 1 0 20944 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_187
timestamp 1669390400
transform 1 0 22288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_194
timestamp 1669390400
transform 1 0 23072 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_196
timestamp 1669390400
transform 1 0 23296 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_205
timestamp 1669390400
transform 1 0 24304 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_224
timestamp 1669390400
transform 1 0 26432 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_234
timestamp 1669390400
transform 1 0 27552 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_244
timestamp 1669390400
transform 1 0 28672 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_246
timestamp 1669390400
transform 1 0 28896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_276
timestamp 1669390400
transform 1 0 32256 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_296
timestamp 1669390400
transform 1 0 34496 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_302
timestamp 1669390400
transform 1 0 35168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_306
timestamp 1669390400
transform 1 0 35616 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_312
timestamp 1669390400
transform 1 0 36288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_326
timestamp 1669390400
transform 1 0 37856 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_333
timestamp 1669390400
transform 1 0 38640 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_343
timestamp 1669390400
transform 1 0 39760 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_347
timestamp 1669390400
transform 1 0 40208 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_363
timestamp 1669390400
transform 1 0 42000 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_365
timestamp 1669390400
transform 1 0 42224 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_69
timestamp 1669390400
transform 1 0 9072 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_72
timestamp 1669390400
transform 1 0 9408 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_76
timestamp 1669390400
transform 1 0 9856 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_80
timestamp 1669390400
transform 1 0 10304 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_84
timestamp 1669390400
transform 1 0 10752 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_88
timestamp 1669390400
transform 1 0 11200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_92
timestamp 1669390400
transform 1 0 11648 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_96
timestamp 1669390400
transform 1 0 12096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_100
timestamp 1669390400
transform 1 0 12544 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_102
timestamp 1669390400
transform 1 0 12768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_111
timestamp 1669390400
transform 1 0 13776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_115
timestamp 1669390400
transform 1 0 14224 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_119
timestamp 1669390400
transform 1 0 14672 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_123
timestamp 1669390400
transform 1 0 15120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_129
timestamp 1669390400
transform 1 0 15792 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_133
timestamp 1669390400
transform 1 0 16240 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_137
timestamp 1669390400
transform 1 0 16688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_141
timestamp 1669390400
transform 1 0 17136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_145
timestamp 1669390400
transform 1 0 17584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_149
timestamp 1669390400
transform 1 0 18032 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_152
timestamp 1669390400
transform 1 0 18368 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_156
timestamp 1669390400
transform 1 0 18816 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_160
timestamp 1669390400
transform 1 0 19264 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_164
timestamp 1669390400
transform 1 0 19712 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_171
timestamp 1669390400
transform 1 0 20496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_173
timestamp 1669390400
transform 1 0 20720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_209
timestamp 1669390400
transform 1 0 24752 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_217
timestamp 1669390400
transform 1 0 25648 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_221
timestamp 1669390400
transform 1 0 26096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_227
timestamp 1669390400
transform 1 0 26768 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_234
timestamp 1669390400
transform 1 0 27552 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_238
timestamp 1669390400
transform 1 0 28000 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_240
timestamp 1669390400
transform 1 0 28224 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_256
timestamp 1669390400
transform 1 0 30016 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_263
timestamp 1669390400
transform 1 0 30800 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_270
timestamp 1669390400
transform 1 0 31584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_283
timestamp 1669390400
transform 1 0 33040 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_290
timestamp 1669390400
transform 1 0 33824 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_296
timestamp 1669390400
transform 1 0 34496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_302
timestamp 1669390400
transform 1 0 35168 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_306
timestamp 1669390400
transform 1 0 35616 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_308
timestamp 1669390400
transform 1 0 35840 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_316
timestamp 1669390400
transform 1 0 36736 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_326
timestamp 1669390400
transform 1 0 37856 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_330
timestamp 1669390400
transform 1 0 38304 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_332
timestamp 1669390400
transform 1 0 38528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_338
timestamp 1669390400
transform 1 0 39200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1669390400
transform 1 0 40096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_353
timestamp 1669390400
transform 1 0 40880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_357
timestamp 1669390400
transform 1 0 41328 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_363
timestamp 1669390400
transform 1 0 42000 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_365
timestamp 1669390400
transform 1 0 42224 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_89
timestamp 1669390400
transform 1 0 11312 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_93
timestamp 1669390400
transform 1 0 11760 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_97
timestamp 1669390400
transform 1 0 12208 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_101
timestamp 1669390400
transform 1 0 12656 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_105
timestamp 1669390400
transform 1 0 13104 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_109
timestamp 1669390400
transform 1 0 13552 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_113
timestamp 1669390400
transform 1 0 14000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_117
timestamp 1669390400
transform 1 0 14448 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_120
timestamp 1669390400
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_126
timestamp 1669390400
transform 1 0 15456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_130
timestamp 1669390400
transform 1 0 15904 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_134
timestamp 1669390400
transform 1 0 16352 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_146
timestamp 1669390400
transform 1 0 17696 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_149
timestamp 1669390400
transform 1 0 18032 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_153
timestamp 1669390400
transform 1 0 18480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_157
timestamp 1669390400
transform 1 0 18928 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_161
timestamp 1669390400
transform 1 0 19376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_165
timestamp 1669390400
transform 1 0 19824 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_168
timestamp 1669390400
transform 1 0 20160 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_199
timestamp 1669390400
transform 1 0 23632 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_206
timestamp 1669390400
transform 1 0 24416 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_210
timestamp 1669390400
transform 1 0 24864 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_224
timestamp 1669390400
transform 1 0 26432 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_226
timestamp 1669390400
transform 1 0 26656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_234
timestamp 1669390400
transform 1 0 27552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_238
timestamp 1669390400
transform 1 0 28000 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_246
timestamp 1669390400
transform 1 0 28896 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_257
timestamp 1669390400
transform 1 0 30128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_264
timestamp 1669390400
transform 1 0 30912 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_266
timestamp 1669390400
transform 1 0 31136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_273
timestamp 1669390400
transform 1 0 31920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_280
timestamp 1669390400
transform 1 0 32704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_292
timestamp 1669390400
transform 1 0 34048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_302
timestamp 1669390400
transform 1 0 35168 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_309
timestamp 1669390400
transform 1 0 35952 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_316
timestamp 1669390400
transform 1 0 36736 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_323
timestamp 1669390400
transform 1 0 37520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_327
timestamp 1669390400
transform 1 0 37968 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_337
timestamp 1669390400
transform 1 0 39088 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_344
timestamp 1669390400
transform 1 0 39872 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_351
timestamp 1669390400
transform 1 0 40656 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_364
timestamp 1669390400
transform 1 0 42112 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_118
timestamp 1669390400
transform 1 0 14560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_122
timestamp 1669390400
transform 1 0 15008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_126
timestamp 1669390400
transform 1 0 15456 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_130
timestamp 1669390400
transform 1 0 15904 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_134
timestamp 1669390400
transform 1 0 16352 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_138
timestamp 1669390400
transform 1 0 16800 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_142
timestamp 1669390400
transform 1 0 17248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_146
timestamp 1669390400
transform 1 0 17696 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_150
timestamp 1669390400
transform 1 0 18144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_154
timestamp 1669390400
transform 1 0 18592 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_157
timestamp 1669390400
transform 1 0 18928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_161
timestamp 1669390400
transform 1 0 19376 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_165
timestamp 1669390400
transform 1 0 19824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_169
timestamp 1669390400
transform 1 0 20272 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_188
timestamp 1669390400
transform 1 0 22400 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_190
timestamp 1669390400
transform 1 0 22624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_200
timestamp 1669390400
transform 1 0 23744 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_210
timestamp 1669390400
transform 1 0 24864 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_221
timestamp 1669390400
transform 1 0 26096 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_225
timestamp 1669390400
transform 1 0 26544 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_235
timestamp 1669390400
transform 1 0 27664 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_246
timestamp 1669390400
transform 1 0 28896 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_258
timestamp 1669390400
transform 1 0 30240 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_264
timestamp 1669390400
transform 1 0 30912 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_274
timestamp 1669390400
transform 1 0 32032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_287
timestamp 1669390400
transform 1 0 33488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_293
timestamp 1669390400
transform 1 0 34160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_300
timestamp 1669390400
transform 1 0 34944 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_307
timestamp 1669390400
transform 1 0 35728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_316
timestamp 1669390400
transform 1 0 36736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_329
timestamp 1669390400
transform 1 0 38192 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_338
timestamp 1669390400
transform 1 0 39200 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_346
timestamp 1669390400
transform 1 0 40096 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_352
timestamp 1669390400
transform 1 0 40768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_356
timestamp 1669390400
transform 1 0 41216 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_363
timestamp 1669390400
transform 1 0 42000 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_365
timestamp 1669390400
transform 1 0 42224 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_105
timestamp 1669390400
transform 1 0 13104 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_121
timestamp 1669390400
transform 1 0 14896 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_125
timestamp 1669390400
transform 1 0 15344 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_147
timestamp 1669390400
transform 1 0 17808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_149
timestamp 1669390400
transform 1 0 18032 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_152
timestamp 1669390400
transform 1 0 18368 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_156
timestamp 1669390400
transform 1 0 18816 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_160
timestamp 1669390400
transform 1 0 19264 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_164
timestamp 1669390400
transform 1 0 19712 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_168
timestamp 1669390400
transform 1 0 20160 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_172
timestamp 1669390400
transform 1 0 20608 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_176
timestamp 1669390400
transform 1 0 21056 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_180
timestamp 1669390400
transform 1 0 21504 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_184
timestamp 1669390400
transform 1 0 21952 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_188
timestamp 1669390400
transform 1 0 22400 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_192
timestamp 1669390400
transform 1 0 22848 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_199
timestamp 1669390400
transform 1 0 23632 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_201
timestamp 1669390400
transform 1 0 23856 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_207
timestamp 1669390400
transform 1 0 24528 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_209
timestamp 1669390400
transform 1 0 24752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_224
timestamp 1669390400
transform 1 0 26432 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_257
timestamp 1669390400
transform 1 0 30128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_266
timestamp 1669390400
transform 1 0 31136 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_273
timestamp 1669390400
transform 1 0 31920 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_280
timestamp 1669390400
transform 1 0 32704 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_316
timestamp 1669390400
transform 1 0 36736 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_326
timestamp 1669390400
transform 1 0 37856 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_328
timestamp 1669390400
transform 1 0 38080 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_337
timestamp 1669390400
transform 1 0 39088 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_344
timestamp 1669390400
transform 1 0 39872 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_352
timestamp 1669390400
transform 1 0 40768 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_364
timestamp 1669390400
transform 1 0 42112 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_140
timestamp 1669390400
transform 1 0 17024 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_148
timestamp 1669390400
transform 1 0 17920 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_152
timestamp 1669390400
transform 1 0 18368 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_155
timestamp 1669390400
transform 1 0 18704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_159
timestamp 1669390400
transform 1 0 19152 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_163
timestamp 1669390400
transform 1 0 19600 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_167
timestamp 1669390400
transform 1 0 20048 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_171
timestamp 1669390400
transform 1 0 20496 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_173
timestamp 1669390400
transform 1 0 20720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_188
timestamp 1669390400
transform 1 0 22400 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_192
timestamp 1669390400
transform 1 0 22848 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_195
timestamp 1669390400
transform 1 0 23184 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_204
timestamp 1669390400
transform 1 0 24192 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_206
timestamp 1669390400
transform 1 0 24416 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_212
timestamp 1669390400
transform 1 0 25088 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_222
timestamp 1669390400
transform 1 0 26208 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_229
timestamp 1669390400
transform 1 0 26992 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_235
timestamp 1669390400
transform 1 0 27664 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_241
timestamp 1669390400
transform 1 0 28336 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_245
timestamp 1669390400
transform 1 0 28784 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_260
timestamp 1669390400
transform 1 0 30464 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_270
timestamp 1669390400
transform 1 0 31584 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_274
timestamp 1669390400
transform 1 0 32032 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_305
timestamp 1669390400
transform 1 0 35504 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_307
timestamp 1669390400
transform 1 0 35728 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_313
timestamp 1669390400
transform 1 0 36400 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_317
timestamp 1669390400
transform 1 0 36848 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_326
timestamp 1669390400
transform 1 0 37856 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_335
timestamp 1669390400
transform 1 0 38864 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_341
timestamp 1669390400
transform 1 0 39536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_347
timestamp 1669390400
transform 1 0 40208 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_353
timestamp 1669390400
transform 1 0 40880 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_359
timestamp 1669390400
transform 1 0 41552 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_365
timestamp 1669390400
transform 1 0 42224 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_160
timestamp 1669390400
transform 1 0 19264 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_164
timestamp 1669390400
transform 1 0 19712 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_168
timestamp 1669390400
transform 1 0 20160 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_199
timestamp 1669390400
transform 1 0 23632 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_209
timestamp 1669390400
transform 1 0 24752 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_248
timestamp 1669390400
transform 1 0 29120 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_257
timestamp 1669390400
transform 1 0 30128 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_263
timestamp 1669390400
transform 1 0 30800 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_267
timestamp 1669390400
transform 1 0 31248 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_271
timestamp 1669390400
transform 1 0 31696 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_275
timestamp 1669390400
transform 1 0 32144 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_289
timestamp 1669390400
transform 1 0 33712 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_293
timestamp 1669390400
transform 1 0 34160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_297
timestamp 1669390400
transform 1 0 34608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_302
timestamp 1669390400
transform 1 0 35168 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_306
timestamp 1669390400
transform 1 0 35616 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_310
timestamp 1669390400
transform 1 0 36064 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_316
timestamp 1669390400
transform 1 0 36736 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_322
timestamp 1669390400
transform 1 0 37408 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_326
timestamp 1669390400
transform 1 0 37856 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_330
timestamp 1669390400
transform 1 0 38304 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_334
timestamp 1669390400
transform 1 0 38752 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_338
timestamp 1669390400
transform 1 0 39200 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_342
timestamp 1669390400
transform 1 0 39648 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_346
timestamp 1669390400
transform 1 0 40096 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_365
timestamp 1669390400
transform 1 0 42224 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_182
timestamp 1669390400
transform 1 0 21728 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_186
timestamp 1669390400
transform 1 0 22176 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_190
timestamp 1669390400
transform 1 0 22624 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_194
timestamp 1669390400
transform 1 0 23072 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_201
timestamp 1669390400
transform 1 0 23856 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_205
timestamp 1669390400
transform 1 0 24304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_209
timestamp 1669390400
transform 1 0 24752 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_217
timestamp 1669390400
transform 1 0 25648 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_224
timestamp 1669390400
transform 1 0 26432 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_228
timestamp 1669390400
transform 1 0 26880 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_232
timestamp 1669390400
transform 1 0 27328 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_234
timestamp 1669390400
transform 1 0 27552 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_237
timestamp 1669390400
transform 1 0 27888 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_241
timestamp 1669390400
transform 1 0 28336 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_245
timestamp 1669390400
transform 1 0 28784 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_253
timestamp 1669390400
transform 1 0 29680 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_257
timestamp 1669390400
transform 1 0 30128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_261
timestamp 1669390400
transform 1 0 30576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_264
timestamp 1669390400
transform 1 0 30912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_268
timestamp 1669390400
transform 1 0 31360 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_272
timestamp 1669390400
transform 1 0 31808 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_278
timestamp 1669390400
transform 1 0 32480 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_282
timestamp 1669390400
transform 1 0 32928 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_286
timestamp 1669390400
transform 1 0 33376 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_290
timestamp 1669390400
transform 1 0 33824 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_292
timestamp 1669390400
transform 1 0 34048 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_295
timestamp 1669390400
transform 1 0 34384 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_299
timestamp 1669390400
transform 1 0 34832 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_303
timestamp 1669390400
transform 1 0 35280 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_309
timestamp 1669390400
transform 1 0 35952 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_313
timestamp 1669390400
transform 1 0 36400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_317
timestamp 1669390400
transform 1 0 36848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_324
timestamp 1669390400
transform 1 0 37632 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_328
timestamp 1669390400
transform 1 0 38080 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_332
timestamp 1669390400
transform 1 0 38528 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_336
timestamp 1669390400
transform 1 0 38976 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_340
timestamp 1669390400
transform 1 0 39424 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_344
timestamp 1669390400
transform 1 0 39872 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_346
timestamp 1669390400
transform 1 0 40096 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_349
timestamp 1669390400
transform 1 0 40432 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_353
timestamp 1669390400
transform 1 0 40880 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_357
timestamp 1669390400
transform 1 0 41328 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_361
timestamp 1669390400
transform 1 0 41776 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_365
timestamp 1669390400
transform 1 0 42224 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_176
timestamp 1669390400
transform 1 0 21056 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_186
timestamp 1669390400
transform 1 0 22176 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_190
timestamp 1669390400
transform 1 0 22624 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_194
timestamp 1669390400
transform 1 0 23072 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_198
timestamp 1669390400
transform 1 0 23520 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_202
timestamp 1669390400
transform 1 0 23968 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_206
timestamp 1669390400
transform 1 0 24416 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_210
timestamp 1669390400
transform 1 0 24864 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_218
timestamp 1669390400
transform 1 0 25760 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_222
timestamp 1669390400
transform 1 0 26208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_226
timestamp 1669390400
transform 1 0 26656 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_230
timestamp 1669390400
transform 1 0 27104 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_234
timestamp 1669390400
transform 1 0 27552 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_238
timestamp 1669390400
transform 1 0 28000 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_242
timestamp 1669390400
transform 1 0 28448 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_246
timestamp 1669390400
transform 1 0 28896 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_250
timestamp 1669390400
transform 1 0 29344 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_254
timestamp 1669390400
transform 1 0 29792 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_258
timestamp 1669390400
transform 1 0 30240 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_262
timestamp 1669390400
transform 1 0 30688 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_266
timestamp 1669390400
transform 1 0 31136 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_270
timestamp 1669390400
transform 1 0 31584 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_274
timestamp 1669390400
transform 1 0 32032 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_278
timestamp 1669390400
transform 1 0 32480 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_282
timestamp 1669390400
transform 1 0 32928 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_289
timestamp 1669390400
transform 1 0 33712 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_293
timestamp 1669390400
transform 1 0 34160 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_297
timestamp 1669390400
transform 1 0 34608 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_301
timestamp 1669390400
transform 1 0 35056 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_305
timestamp 1669390400
transform 1 0 35504 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_309
timestamp 1669390400
transform 1 0 35952 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_313
timestamp 1669390400
transform 1 0 36400 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_317
timestamp 1669390400
transform 1 0 36848 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_321
timestamp 1669390400
transform 1 0 37296 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_325
timestamp 1669390400
transform 1 0 37744 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_329
timestamp 1669390400
transform 1 0 38192 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_333
timestamp 1669390400
transform 1 0 38640 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_337
timestamp 1669390400
transform 1 0 39088 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_341
timestamp 1669390400
transform 1 0 39536 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_345
timestamp 1669390400
transform 1 0 39984 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_347
timestamp 1669390400
transform 1 0 40208 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_360
timestamp 1669390400
transform 1 0 41664 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_364
timestamp 1669390400
transform 1 0 42112 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_187
timestamp 1669390400
transform 1 0 22288 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_191
timestamp 1669390400
transform 1 0 22736 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_194
timestamp 1669390400
transform 1 0 23072 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_198
timestamp 1669390400
transform 1 0 23520 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_202
timestamp 1669390400
transform 1 0 23968 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_206
timestamp 1669390400
transform 1 0 24416 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_210
timestamp 1669390400
transform 1 0 24864 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_214
timestamp 1669390400
transform 1 0 25312 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_216
timestamp 1669390400
transform 1 0 25536 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_219
timestamp 1669390400
transform 1 0 25872 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_223
timestamp 1669390400
transform 1 0 26320 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_227
timestamp 1669390400
transform 1 0 26768 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_231
timestamp 1669390400
transform 1 0 27216 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_235
timestamp 1669390400
transform 1 0 27664 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_238
timestamp 1669390400
transform 1 0 28000 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_242
timestamp 1669390400
transform 1 0 28448 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1669390400
transform 1 0 28896 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_253
timestamp 1669390400
transform 1 0 29680 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_257
timestamp 1669390400
transform 1 0 30128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_261
timestamp 1669390400
transform 1 0 30576 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_265
timestamp 1669390400
transform 1 0 31024 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_269
timestamp 1669390400
transform 1 0 31472 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_273
timestamp 1669390400
transform 1 0 31920 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_277
timestamp 1669390400
transform 1 0 32368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_281
timestamp 1669390400
transform 1 0 32816 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_285
timestamp 1669390400
transform 1 0 33264 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_289
timestamp 1669390400
transform 1 0 33712 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_293
timestamp 1669390400
transform 1 0 34160 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_297
timestamp 1669390400
transform 1 0 34608 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_301
timestamp 1669390400
transform 1 0 35056 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_305
timestamp 1669390400
transform 1 0 35504 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_309
timestamp 1669390400
transform 1 0 35952 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_313
timestamp 1669390400
transform 1 0 36400 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1669390400
transform 1 0 36848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_324
timestamp 1669390400
transform 1 0 37632 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_328
timestamp 1669390400
transform 1 0 38080 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_332
timestamp 1669390400
transform 1 0 38528 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_336
timestamp 1669390400
transform 1 0 38976 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_340
timestamp 1669390400
transform 1 0 39424 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_344
timestamp 1669390400
transform 1 0 39872 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_347
timestamp 1669390400
transform 1 0 40208 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_351
timestamp 1669390400
transform 1 0 40656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_355
timestamp 1669390400
transform 1 0 41104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_358
timestamp 1669390400
transform 1 0 41440 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_362
timestamp 1669390400
transform 1 0 41888 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_365
timestamp 1669390400
transform 1 0 42224 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_5
timestamp 1669390400
transform 1 0 1904 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_69
timestamp 1669390400
transform 1 0 9072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_176
timestamp 1669390400
transform 1 0 21056 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_192
timestamp 1669390400
transform 1 0 22848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_200
timestamp 1669390400
transform 1 0 23744 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_204
timestamp 1669390400
transform 1 0 24192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_218
timestamp 1669390400
transform 1 0 25760 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_220
timestamp 1669390400
transform 1 0 25984 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_223
timestamp 1669390400
transform 1 0 26320 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_227
timestamp 1669390400
transform 1 0 26768 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_231
timestamp 1669390400
transform 1 0 27216 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_235
timestamp 1669390400
transform 1 0 27664 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_239
timestamp 1669390400
transform 1 0 28112 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_243
timestamp 1669390400
transform 1 0 28560 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_247
timestamp 1669390400
transform 1 0 29008 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_251
timestamp 1669390400
transform 1 0 29456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_255
timestamp 1669390400
transform 1 0 29904 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_258
timestamp 1669390400
transform 1 0 30240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_262
timestamp 1669390400
transform 1 0 30688 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_266
timestamp 1669390400
transform 1 0 31136 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_270
timestamp 1669390400
transform 1 0 31584 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_273
timestamp 1669390400
transform 1 0 31920 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_277
timestamp 1669390400
transform 1 0 32368 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_281
timestamp 1669390400
transform 1 0 32816 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_289
timestamp 1669390400
transform 1 0 33712 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_293
timestamp 1669390400
transform 1 0 34160 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_297
timestamp 1669390400
transform 1 0 34608 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_301
timestamp 1669390400
transform 1 0 35056 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_305
timestamp 1669390400
transform 1 0 35504 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_309
timestamp 1669390400
transform 1 0 35952 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_313
timestamp 1669390400
transform 1 0 36400 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_317
timestamp 1669390400
transform 1 0 36848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_321
timestamp 1669390400
transform 1 0 37296 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_325
timestamp 1669390400
transform 1 0 37744 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_329
timestamp 1669390400
transform 1 0 38192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_333
timestamp 1669390400
transform 1 0 38640 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_337
timestamp 1669390400
transform 1 0 39088 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_341
timestamp 1669390400
transform 1 0 39536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_347
timestamp 1669390400
transform 1 0 40208 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_351
timestamp 1669390400
transform 1 0 40656 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_360
timestamp 1669390400
transform 1 0 41664 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_362
timestamp 1669390400
transform 1 0 41888 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_365
timestamp 1669390400
transform 1 0 42224 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_19
timestamp 1669390400
transform 1 0 3472 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_195
timestamp 1669390400
transform 1 0 23184 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_203
timestamp 1669390400
transform 1 0 24080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_207
timestamp 1669390400
transform 1 0 24528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_210
timestamp 1669390400
transform 1 0 24864 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_214
timestamp 1669390400
transform 1 0 25312 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_218
timestamp 1669390400
transform 1 0 25760 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_222
timestamp 1669390400
transform 1 0 26208 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_226
timestamp 1669390400
transform 1 0 26656 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_230
timestamp 1669390400
transform 1 0 27104 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_234
timestamp 1669390400
transform 1 0 27552 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_238
timestamp 1669390400
transform 1 0 28000 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_244
timestamp 1669390400
transform 1 0 28672 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_253
timestamp 1669390400
transform 1 0 29680 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_257
timestamp 1669390400
transform 1 0 30128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_261
timestamp 1669390400
transform 1 0 30576 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_265
timestamp 1669390400
transform 1 0 31024 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_269
timestamp 1669390400
transform 1 0 31472 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_273
timestamp 1669390400
transform 1 0 31920 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_277
timestamp 1669390400
transform 1 0 32368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_281
timestamp 1669390400
transform 1 0 32816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_287
timestamp 1669390400
transform 1 0 33488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_291
timestamp 1669390400
transform 1 0 33936 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_295
timestamp 1669390400
transform 1 0 34384 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_299
timestamp 1669390400
transform 1 0 34832 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_303
timestamp 1669390400
transform 1 0 35280 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_307
timestamp 1669390400
transform 1 0 35728 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_311
timestamp 1669390400
transform 1 0 36176 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_315
timestamp 1669390400
transform 1 0 36624 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_324
timestamp 1669390400
transform 1 0 37632 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_328
timestamp 1669390400
transform 1 0 38080 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_332
timestamp 1669390400
transform 1 0 38528 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_348
timestamp 1669390400
transform 1 0 40320 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_352
timestamp 1669390400
transform 1 0 40768 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_356
timestamp 1669390400
transform 1 0 41216 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_358
timestamp 1669390400
transform 1 0 41440 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_361
timestamp 1669390400
transform 1 0 41776 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_365
timestamp 1669390400
transform 1 0 42224 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_219
timestamp 1669390400
transform 1 0 25872 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_223
timestamp 1669390400
transform 1 0 26320 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_227
timestamp 1669390400
transform 1 0 26768 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_231
timestamp 1669390400
transform 1 0 27216 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_235
timestamp 1669390400
transform 1 0 27664 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_241
timestamp 1669390400
transform 1 0 28336 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_245
timestamp 1669390400
transform 1 0 28784 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_251
timestamp 1669390400
transform 1 0 29456 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_255
timestamp 1669390400
transform 1 0 29904 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_261
timestamp 1669390400
transform 1 0 30576 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_265
timestamp 1669390400
transform 1 0 31024 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_271
timestamp 1669390400
transform 1 0 31696 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_275
timestamp 1669390400
transform 1 0 32144 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_289
timestamp 1669390400
transform 1 0 33712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_293
timestamp 1669390400
transform 1 0 34160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_297
timestamp 1669390400
transform 1 0 34608 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_301
timestamp 1669390400
transform 1 0 35056 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_305
timestamp 1669390400
transform 1 0 35504 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_309
timestamp 1669390400
transform 1 0 35952 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_313
timestamp 1669390400
transform 1 0 36400 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_317
timestamp 1669390400
transform 1 0 36848 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_321
timestamp 1669390400
transform 1 0 37296 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_325
timestamp 1669390400
transform 1 0 37744 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_331
timestamp 1669390400
transform 1 0 38416 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_335
timestamp 1669390400
transform 1 0 38864 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_337
timestamp 1669390400
transform 1 0 39088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_340
timestamp 1669390400
transform 1 0 39424 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_344
timestamp 1669390400
transform 1 0 39872 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_348
timestamp 1669390400
transform 1 0 40320 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_352
timestamp 1669390400
transform 1 0 40768 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_360
timestamp 1669390400
transform 1 0 41664 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_362
timestamp 1669390400
transform 1 0 41888 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_365
timestamp 1669390400
transform 1 0 42224 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_211
timestamp 1669390400
transform 1 0 24976 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_227
timestamp 1669390400
transform 1 0 26768 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_235
timestamp 1669390400
transform 1 0 27664 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_239
timestamp 1669390400
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_245
timestamp 1669390400
transform 1 0 28784 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_253
timestamp 1669390400
transform 1 0 29680 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_257
timestamp 1669390400
transform 1 0 30128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_261
timestamp 1669390400
transform 1 0 30576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_267
timestamp 1669390400
transform 1 0 31248 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_271
timestamp 1669390400
transform 1 0 31696 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_275
timestamp 1669390400
transform 1 0 32144 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_279
timestamp 1669390400
transform 1 0 32592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_283
timestamp 1669390400
transform 1 0 33040 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_287
timestamp 1669390400
transform 1 0 33488 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_291
timestamp 1669390400
transform 1 0 33936 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_295
timestamp 1669390400
transform 1 0 34384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_299
timestamp 1669390400
transform 1 0 34832 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_301
timestamp 1669390400
transform 1 0 35056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_304
timestamp 1669390400
transform 1 0 35392 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_308
timestamp 1669390400
transform 1 0 35840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_323
timestamp 1669390400
transform 1 0 37520 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_326
timestamp 1669390400
transform 1 0 37856 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_330
timestamp 1669390400
transform 1 0 38304 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_334
timestamp 1669390400
transform 1 0 38752 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_338
timestamp 1669390400
transform 1 0 39200 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_342
timestamp 1669390400
transform 1 0 39648 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_348
timestamp 1669390400
transform 1 0 40320 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_352
timestamp 1669390400
transform 1 0 40768 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_358
timestamp 1669390400
transform 1 0 41440 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_362
timestamp 1669390400
transform 1 0 41888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_247
timestamp 1669390400
transform 1 0 29008 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_255
timestamp 1669390400
transform 1 0 29904 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_258
timestamp 1669390400
transform 1 0 30240 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_262
timestamp 1669390400
transform 1 0 30688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_270
timestamp 1669390400
transform 1 0 31584 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_273
timestamp 1669390400
transform 1 0 31920 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_281
timestamp 1669390400
transform 1 0 32816 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_360
timestamp 1669390400
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_364
timestamp 1669390400
transform 1 0 42112 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_353
timestamp 1669390400
transform 1 0 40880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_361
timestamp 1669390400
transform 1 0 41776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_365
timestamp 1669390400
transform 1 0 42224 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_365
timestamp 1669390400
transform 1 0 42224 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_353
timestamp 1669390400
transform 1 0 40880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_361
timestamp 1669390400
transform 1 0 41776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_365
timestamp 1669390400
transform 1 0 42224 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_365
timestamp 1669390400
transform 1 0 42224 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_353
timestamp 1669390400
transform 1 0 40880 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_361
timestamp 1669390400
transform 1 0 41776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_365
timestamp 1669390400
transform 1 0 42224 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_365
timestamp 1669390400
transform 1 0 42224 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_353
timestamp 1669390400
transform 1 0 40880 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_361
timestamp 1669390400
transform 1 0 41776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_365
timestamp 1669390400
transform 1 0 42224 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_365
timestamp 1669390400
transform 1 0 42224 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_353
timestamp 1669390400
transform 1 0 40880 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_361
timestamp 1669390400
transform 1 0 41776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_365
timestamp 1669390400
transform 1 0 42224 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_365
timestamp 1669390400
transform 1 0 42224 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_353
timestamp 1669390400
transform 1 0 40880 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_361
timestamp 1669390400
transform 1 0 41776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_365
timestamp 1669390400
transform 1 0 42224 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_365
timestamp 1669390400
transform 1 0 42224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_353
timestamp 1669390400
transform 1 0 40880 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_361
timestamp 1669390400
transform 1 0 41776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_365
timestamp 1669390400
transform 1 0 42224 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_365
timestamp 1669390400
transform 1 0 42224 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_353
timestamp 1669390400
transform 1 0 40880 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_361
timestamp 1669390400
transform 1 0 41776 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_365
timestamp 1669390400
transform 1 0 42224 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_365
timestamp 1669390400
transform 1 0 42224 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_353
timestamp 1669390400
transform 1 0 40880 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_361
timestamp 1669390400
transform 1 0 41776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_365
timestamp 1669390400
transform 1 0 42224 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_353
timestamp 1669390400
transform 1 0 40880 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_361
timestamp 1669390400
transform 1 0 41776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_365
timestamp 1669390400
transform 1 0 42224 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_34
timestamp 1669390400
transform 1 0 5152 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_37
timestamp 1669390400
transform 1 0 5488 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_69
timestamp 1669390400
transform 1 0 9072 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_72
timestamp 1669390400
transform 1 0 9408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_104
timestamp 1669390400
transform 1 0 12992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_107
timestamp 1669390400
transform 1 0 13328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_139
timestamp 1669390400
transform 1 0 16912 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_142
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_174
timestamp 1669390400
transform 1 0 20832 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_177
timestamp 1669390400
transform 1 0 21168 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_209
timestamp 1669390400
transform 1 0 24752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_244
timestamp 1669390400
transform 1 0 28672 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_247
timestamp 1669390400
transform 1 0 29008 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_282
timestamp 1669390400
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_314
timestamp 1669390400
transform 1 0 36512 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_317
timestamp 1669390400
transform 1 0 36848 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_349
timestamp 1669390400
transform 1 0 40432 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_352
timestamp 1669390400
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_360
timestamp 1669390400
transform 1 0 41664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_364
timestamp 1669390400
transform 1 0 42112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 42560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 42560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 42560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 42560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 42560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 42560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 42560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 42560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 42560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 42560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 42560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 42560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 42560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 42560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 42560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 42560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 42560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 42560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 42560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 42560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 42560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 42560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 42560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 42560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 42560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 42560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 42560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 42560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 42560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 42560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 42560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 42560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 5264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 13104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 20944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 28784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 36624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _344_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24976 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _345_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 21056 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _346_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30240 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _347_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29456 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _348_
timestamp 1669390400
transform 1 0 15232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _349_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _350_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5936 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _351_
timestamp 1669390400
transform -1 0 36960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _352_
timestamp 1669390400
transform -1 0 30016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _353_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4256 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _354_
timestamp 1669390400
transform -1 0 3360 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _355_
timestamp 1669390400
transform -1 0 6160 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _356_
timestamp 1669390400
transform 1 0 4032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _357_
timestamp 1669390400
transform -1 0 7056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _358_
timestamp 1669390400
transform -1 0 5040 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _359_
timestamp 1669390400
transform 1 0 30688 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _360_
timestamp 1669390400
transform 1 0 31696 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _361_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6496 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _362_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3472 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _363_
timestamp 1669390400
transform -1 0 8512 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _364_
timestamp 1669390400
transform 1 0 4480 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _365_
timestamp 1669390400
transform -1 0 10976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _366_
timestamp 1669390400
transform -1 0 8736 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _367_
timestamp 1669390400
transform -1 0 12992 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _368_
timestamp 1669390400
transform 1 0 4368 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _369_
timestamp 1669390400
transform 1 0 7616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _370_
timestamp 1669390400
transform 1 0 10528 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _371_
timestamp 1669390400
transform -1 0 13104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _372_
timestamp 1669390400
transform 1 0 12432 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _373_
timestamp 1669390400
transform 1 0 13552 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _374_
timestamp 1669390400
transform 1 0 14224 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _375_
timestamp 1669390400
transform -1 0 18032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _376_
timestamp 1669390400
transform 1 0 8960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _377_
timestamp 1669390400
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _378_
timestamp 1669390400
transform -1 0 14336 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _379_
timestamp 1669390400
transform -1 0 18704 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _380_
timestamp 1669390400
transform -1 0 14336 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _381_
timestamp 1669390400
transform -1 0 18480 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _382_
timestamp 1669390400
transform -1 0 18368 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _383_
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _384_
timestamp 1669390400
transform 1 0 19488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _385_
timestamp 1669390400
transform -1 0 24304 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _386_
timestamp 1669390400
transform -1 0 37632 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _387_
timestamp 1669390400
transform -1 0 22400 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _388_
timestamp 1669390400
transform 1 0 19936 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _389_
timestamp 1669390400
transform 1 0 27776 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _390_
timestamp 1669390400
transform 1 0 21840 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _391_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22736 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _392_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21168 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _393_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 35504 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _394_
timestamp 1669390400
transform -1 0 33040 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _395_
timestamp 1669390400
transform -1 0 42112 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _396_
timestamp 1669390400
transform -1 0 36176 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _397_
timestamp 1669390400
transform -1 0 24528 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _398_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23856 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _399_
timestamp 1669390400
transform 1 0 18704 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _400_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21840 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _401_
timestamp 1669390400
transform -1 0 42112 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _402_
timestamp 1669390400
transform 1 0 40432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _403_
timestamp 1669390400
transform 1 0 41552 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _404_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23968 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _405_
timestamp 1669390400
transform 1 0 35840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _406_
timestamp 1669390400
transform 1 0 36176 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _407_
timestamp 1669390400
transform -1 0 40768 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _408_
timestamp 1669390400
transform -1 0 30912 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _409_
timestamp 1669390400
transform -1 0 30800 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _410_
timestamp 1669390400
transform 1 0 29456 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _411_
timestamp 1669390400
transform 1 0 30352 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _412_
timestamp 1669390400
transform 1 0 23296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _413_
timestamp 1669390400
transform -1 0 30128 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _414_
timestamp 1669390400
transform -1 0 34496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _415_
timestamp 1669390400
transform -1 0 35168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1669390400
transform -1 0 32704 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _417_
timestamp 1669390400
transform 1 0 26320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _418_
timestamp 1669390400
transform 1 0 27552 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _419_
timestamp 1669390400
transform -1 0 35952 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _420_
timestamp 1669390400
transform 1 0 36960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _421_
timestamp 1669390400
transform 1 0 20384 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _422_
timestamp 1669390400
transform -1 0 22624 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _423_
timestamp 1669390400
transform 1 0 20496 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _424_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 35168 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _425_
timestamp 1669390400
transform -1 0 37856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _426_
timestamp 1669390400
transform -1 0 33040 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _427_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 27776 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _428_
timestamp 1669390400
transform -1 0 21056 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _429_
timestamp 1669390400
transform 1 0 27216 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _430_
timestamp 1669390400
transform -1 0 26880 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _431_
timestamp 1669390400
transform -1 0 23072 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _432_
timestamp 1669390400
transform 1 0 14112 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _433_
timestamp 1669390400
transform -1 0 15456 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _434_
timestamp 1669390400
transform -1 0 6160 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _435_
timestamp 1669390400
transform 1 0 4816 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _436_
timestamp 1669390400
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _437_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7168 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _438_
timestamp 1669390400
transform 1 0 3472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _439_
timestamp 1669390400
transform -1 0 7056 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _440_
timestamp 1669390400
transform -1 0 5600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _441_
timestamp 1669390400
transform 1 0 4592 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _442_
timestamp 1669390400
transform -1 0 7392 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _443_
timestamp 1669390400
transform 1 0 5824 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _444_
timestamp 1669390400
transform 1 0 8176 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _445_
timestamp 1669390400
transform 1 0 7280 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _446_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8288 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _447_
timestamp 1669390400
transform 1 0 7504 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _448_
timestamp 1669390400
transform -1 0 9184 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _449_
timestamp 1669390400
transform 1 0 5936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _450_
timestamp 1669390400
transform 1 0 6608 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _451_
timestamp 1669390400
transform 1 0 9520 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _452_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 25088 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _453_
timestamp 1669390400
transform 1 0 27216 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _454_
timestamp 1669390400
transform 1 0 6608 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _455_
timestamp 1669390400
transform 1 0 8512 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _456_
timestamp 1669390400
transform -1 0 11312 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _457_
timestamp 1669390400
transform -1 0 10640 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _458_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10640 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _459_
timestamp 1669390400
transform 1 0 11536 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _460_
timestamp 1669390400
transform 1 0 10752 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _461_
timestamp 1669390400
transform 1 0 11872 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _462_
timestamp 1669390400
transform -1 0 12320 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _463_
timestamp 1669390400
transform 1 0 7280 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _464_
timestamp 1669390400
transform -1 0 13104 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _465_
timestamp 1669390400
transform 1 0 11088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _466_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 12096 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _467_
timestamp 1669390400
transform 1 0 5600 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _468_
timestamp 1669390400
transform -1 0 11872 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _469_
timestamp 1669390400
transform 1 0 11760 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _470_
timestamp 1669390400
transform 1 0 10640 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _471_
timestamp 1669390400
transform 1 0 13552 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _472_
timestamp 1669390400
transform -1 0 9184 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _473_
timestamp 1669390400
transform -1 0 10192 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _474_
timestamp 1669390400
transform 1 0 4144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _475_
timestamp 1669390400
transform -1 0 10976 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _476_
timestamp 1669390400
transform 1 0 14560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _477_
timestamp 1669390400
transform 1 0 14896 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _478_
timestamp 1669390400
transform 1 0 15344 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _479_
timestamp 1669390400
transform 1 0 14336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _480_
timestamp 1669390400
transform -1 0 10304 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _481_
timestamp 1669390400
transform -1 0 18032 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _482_
timestamp 1669390400
transform 1 0 13328 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _483_
timestamp 1669390400
transform 1 0 15456 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _484_
timestamp 1669390400
transform -1 0 19936 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _485_
timestamp 1669390400
transform -1 0 10752 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _486_
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _487_
timestamp 1669390400
transform 1 0 19376 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _488_
timestamp 1669390400
transform 1 0 19376 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _489_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17696 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _490_
timestamp 1669390400
transform 1 0 18256 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _491_
timestamp 1669390400
transform 1 0 16464 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _492_
timestamp 1669390400
transform 1 0 19824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _493_
timestamp 1669390400
transform -1 0 19264 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _494_
timestamp 1669390400
transform 1 0 16240 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _495_
timestamp 1669390400
transform -1 0 18704 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _496_
timestamp 1669390400
transform -1 0 19824 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _497_
timestamp 1669390400
transform -1 0 17920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _498_
timestamp 1669390400
transform 1 0 26656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _499_
timestamp 1669390400
transform 1 0 25536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _500_
timestamp 1669390400
transform -1 0 25088 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _501_
timestamp 1669390400
transform 1 0 20160 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _502_
timestamp 1669390400
transform 1 0 23968 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _503_
timestamp 1669390400
transform -1 0 17136 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _504_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21504 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _505_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 24080 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _506_
timestamp 1669390400
transform -1 0 28896 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _507_
timestamp 1669390400
transform -1 0 28112 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _508_
timestamp 1669390400
transform -1 0 31696 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _509_
timestamp 1669390400
transform -1 0 26096 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _510_
timestamp 1669390400
transform -1 0 26992 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _511_
timestamp 1669390400
transform 1 0 24416 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _512_
timestamp 1669390400
transform 1 0 21616 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _513_
timestamp 1669390400
transform 1 0 33488 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _514_
timestamp 1669390400
transform 1 0 18144 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _515_
timestamp 1669390400
transform 1 0 26544 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _516_
timestamp 1669390400
transform -1 0 36288 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _517_
timestamp 1669390400
transform -1 0 26320 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _518_
timestamp 1669390400
transform -1 0 24192 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _519_
timestamp 1669390400
transform -1 0 24864 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _520_
timestamp 1669390400
transform 1 0 22624 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _521_
timestamp 1669390400
transform -1 0 23856 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _522_
timestamp 1669390400
transform -1 0 24976 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _523_
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _524_
timestamp 1669390400
transform 1 0 24752 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _525_
timestamp 1669390400
transform 1 0 21056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _526_
timestamp 1669390400
transform 1 0 29456 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _527_
timestamp 1669390400
transform 1 0 26096 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _528_
timestamp 1669390400
transform 1 0 32704 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _529_
timestamp 1669390400
transform -1 0 29008 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _530_
timestamp 1669390400
transform -1 0 27216 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _531_
timestamp 1669390400
transform 1 0 24304 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _532_
timestamp 1669390400
transform 1 0 25088 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _533_
timestamp 1669390400
transform -1 0 39200 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _534_
timestamp 1669390400
transform 1 0 30352 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _535_
timestamp 1669390400
transform -1 0 34160 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _536_
timestamp 1669390400
transform 1 0 30352 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _537_
timestamp 1669390400
transform 1 0 28336 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _538_
timestamp 1669390400
transform -1 0 28336 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _539_
timestamp 1669390400
transform 1 0 27776 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _540_
timestamp 1669390400
transform 1 0 27216 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _541_
timestamp 1669390400
transform 1 0 26320 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _542_
timestamp 1669390400
transform 1 0 27440 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _543_
timestamp 1669390400
transform -1 0 28000 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _544_
timestamp 1669390400
transform 1 0 30576 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _545_
timestamp 1669390400
transform 1 0 31808 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _546_
timestamp 1669390400
transform 1 0 31248 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _547_
timestamp 1669390400
transform 1 0 33488 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _548_
timestamp 1669390400
transform 1 0 29904 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _549_
timestamp 1669390400
transform 1 0 35728 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _550_
timestamp 1669390400
transform -1 0 31808 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _551_
timestamp 1669390400
transform 1 0 30464 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _552_
timestamp 1669390400
transform 1 0 34720 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _553_
timestamp 1669390400
transform 1 0 29568 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _554_
timestamp 1669390400
transform -1 0 39984 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _555_
timestamp 1669390400
transform -1 0 37968 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _556_
timestamp 1669390400
transform 1 0 34720 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _557_
timestamp 1669390400
transform -1 0 35056 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _558_
timestamp 1669390400
transform 1 0 31360 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _559_
timestamp 1669390400
transform -1 0 37968 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _560_
timestamp 1669390400
transform 1 0 30688 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _561_
timestamp 1669390400
transform -1 0 32480 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _562_
timestamp 1669390400
transform -1 0 32928 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _563_
timestamp 1669390400
transform -1 0 42224 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _564_
timestamp 1669390400
transform 1 0 30800 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _565_
timestamp 1669390400
transform -1 0 36960 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _566_
timestamp 1669390400
transform 1 0 37856 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _567_
timestamp 1669390400
transform 1 0 29456 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _568_
timestamp 1669390400
transform -1 0 28560 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _569_
timestamp 1669390400
transform -1 0 29008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _570_
timestamp 1669390400
transform -1 0 33824 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _571_
timestamp 1669390400
transform 1 0 28336 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _572_
timestamp 1669390400
transform -1 0 42000 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _573_
timestamp 1669390400
transform -1 0 41216 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _574_
timestamp 1669390400
transform 1 0 40432 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _575_
timestamp 1669390400
transform -1 0 42000 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _576_
timestamp 1669390400
transform -1 0 42000 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _577_
timestamp 1669390400
transform 1 0 39760 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _578_
timestamp 1669390400
transform 1 0 41776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _579_
timestamp 1669390400
transform -1 0 42000 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _580_
timestamp 1669390400
transform -1 0 38528 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _581_
timestamp 1669390400
transform 1 0 31360 0 1 3136
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _582_
timestamp 1669390400
transform -1 0 37968 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _583_
timestamp 1669390400
transform -1 0 42000 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _584_
timestamp 1669390400
transform -1 0 42000 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _585_
timestamp 1669390400
transform -1 0 41552 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _586_
timestamp 1669390400
transform -1 0 41552 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _587_
timestamp 1669390400
transform -1 0 39872 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _588_
timestamp 1669390400
transform -1 0 41776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _589_
timestamp 1669390400
transform -1 0 37184 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _590_
timestamp 1669390400
transform 1 0 35840 0 1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _591_
timestamp 1669390400
transform -1 0 39536 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _592_
timestamp 1669390400
transform 1 0 41440 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _593_
timestamp 1669390400
transform 1 0 39424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _594_
timestamp 1669390400
transform -1 0 42000 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _595_
timestamp 1669390400
transform -1 0 41888 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _596_
timestamp 1669390400
transform 1 0 40768 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _597_
timestamp 1669390400
transform -1 0 39200 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _598_
timestamp 1669390400
transform -1 0 42112 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _599_
timestamp 1669390400
transform -1 0 38640 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _600_
timestamp 1669390400
transform 1 0 34496 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _601_
timestamp 1669390400
transform -1 0 36960 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _602_
timestamp 1669390400
transform -1 0 42000 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _603_
timestamp 1669390400
transform -1 0 41104 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _604_
timestamp 1669390400
transform 1 0 37408 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _605_
timestamp 1669390400
transform -1 0 40768 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _606_
timestamp 1669390400
transform 1 0 38080 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _607_
timestamp 1669390400
transform -1 0 37856 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _608_
timestamp 1669390400
transform -1 0 35504 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _609_
timestamp 1669390400
transform 1 0 31920 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _610_
timestamp 1669390400
transform 1 0 38416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _611_
timestamp 1669390400
transform -1 0 42112 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _612_
timestamp 1669390400
transform 1 0 39424 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _613_
timestamp 1669390400
transform -1 0 42000 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _614_
timestamp 1669390400
transform -1 0 39984 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _615_
timestamp 1669390400
transform 1 0 39312 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _616_
timestamp 1669390400
transform -1 0 42224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _617_
timestamp 1669390400
transform -1 0 38752 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _618_
timestamp 1669390400
transform -1 0 40768 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _619_
timestamp 1669390400
transform -1 0 39424 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _620_
timestamp 1669390400
transform -1 0 40208 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _621_
timestamp 1669390400
transform 1 0 40432 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _622_
timestamp 1669390400
transform -1 0 38864 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _623_
timestamp 1669390400
transform -1 0 36176 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _624_
timestamp 1669390400
transform 1 0 33488 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _625_
timestamp 1669390400
transform -1 0 40768 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _626_
timestamp 1669390400
transform 1 0 37520 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1669390400
transform 1 0 35616 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _628_
timestamp 1669390400
transform -1 0 36960 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _629_
timestamp 1669390400
transform -1 0 37408 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _630_
timestamp 1669390400
transform 1 0 35728 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _631_
timestamp 1669390400
transform 1 0 35952 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _632_
timestamp 1669390400
transform 1 0 34048 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _633_
timestamp 1669390400
transform 1 0 32032 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _634_
timestamp 1669390400
transform 1 0 37968 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _635_
timestamp 1669390400
transform -1 0 39760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _636_
timestamp 1669390400
transform 1 0 37184 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _637_
timestamp 1669390400
transform 1 0 39088 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _638_
timestamp 1669390400
transform 1 0 39312 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1669390400
transform 1 0 35392 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _640_
timestamp 1669390400
transform 1 0 35168 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _641_
timestamp 1669390400
transform 1 0 35840 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _642_
timestamp 1669390400
transform -1 0 40768 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _643_
timestamp 1669390400
transform -1 0 39872 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _644_
timestamp 1669390400
transform -1 0 39200 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _645_
timestamp 1669390400
transform -1 0 38864 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _646_
timestamp 1669390400
transform -1 0 34720 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _647_
timestamp 1669390400
transform 1 0 32480 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _648_
timestamp 1669390400
transform -1 0 39088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _649_
timestamp 1669390400
transform 1 0 36288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _650_
timestamp 1669390400
transform -1 0 34944 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _651_
timestamp 1669390400
transform 1 0 36176 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _652_
timestamp 1669390400
transform 1 0 37408 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _653_
timestamp 1669390400
transform 1 0 36960 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _654_
timestamp 1669390400
transform 1 0 37408 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _655_
timestamp 1669390400
transform 1 0 35952 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _656_
timestamp 1669390400
transform -1 0 30016 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1669390400
transform -1 0 29008 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _658_
timestamp 1669390400
transform 1 0 29456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _659_
timestamp 1669390400
transform 1 0 39424 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _660_
timestamp 1669390400
transform 1 0 38640 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _661_
timestamp 1669390400
transform 1 0 39424 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _662_
timestamp 1669390400
transform -1 0 40992 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _663_
timestamp 1669390400
transform -1 0 39984 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _664_
timestamp 1669390400
transform -1 0 40880 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _665_
timestamp 1669390400
transform 1 0 36960 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _666_
timestamp 1669390400
transform -1 0 39088 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _667_
timestamp 1669390400
transform 1 0 40096 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _668_
timestamp 1669390400
transform -1 0 31920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1669390400
transform -1 0 34048 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _670_
timestamp 1669390400
transform -1 0 30800 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _671_
timestamp 1669390400
transform 1 0 32144 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _672_
timestamp 1669390400
transform -1 0 31584 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _673_
timestamp 1669390400
transform -1 0 34160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _674_
timestamp 1669390400
transform 1 0 31136 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _675_
timestamp 1669390400
transform 1 0 26992 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _676_
timestamp 1669390400
transform 1 0 27888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _677_
timestamp 1669390400
transform 1 0 28112 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _678_
timestamp 1669390400
transform 1 0 27888 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _679_
timestamp 1669390400
transform -1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _680_
timestamp 1669390400
transform -1 0 30912 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _681_
timestamp 1669390400
transform -1 0 31920 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _682_
timestamp 1669390400
transform -1 0 30240 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _683_
timestamp 1669390400
transform -1 0 30128 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _684_
timestamp 1669390400
transform -1 0 30128 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _685_
timestamp 1669390400
transform -1 0 27552 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _686_
timestamp 1669390400
transform 1 0 25088 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _687_
timestamp 1669390400
transform 1 0 25536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _688_
timestamp 1669390400
transform 1 0 30352 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _689_
timestamp 1669390400
transform -1 0 30464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _690_
timestamp 1669390400
transform 1 0 30688 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _691_
timestamp 1669390400
transform 1 0 25536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _692_
timestamp 1669390400
transform -1 0 25088 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _693_
timestamp 1669390400
transform 1 0 26432 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _694_
timestamp 1669390400
transform -1 0 27664 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _695_
timestamp 1669390400
transform -1 0 26208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _696_
timestamp 1669390400
transform -1 0 26432 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _697_
timestamp 1669390400
transform 1 0 24864 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _698_
timestamp 1669390400
transform 1 0 22736 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _699_
timestamp 1669390400
transform -1 0 22400 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _700_
timestamp 1669390400
transform -1 0 24416 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _701_
timestamp 1669390400
transform 1 0 23968 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _702_
timestamp 1669390400
transform -1 0 24192 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _703_
timestamp 1669390400
transform -1 0 23856 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _704_
timestamp 1669390400
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _705_
timestamp 1669390400
transform -1 0 23632 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _706_
timestamp 1669390400
transform 1 0 21504 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _707_ gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16800 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _708_
timestamp 1669390400
transform -1 0 9968 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _709_
timestamp 1669390400
transform -1 0 9632 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _710_
timestamp 1669390400
transform -1 0 9744 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _711_
timestamp 1669390400
transform 1 0 5936 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _712_
timestamp 1669390400
transform -1 0 10304 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _713_
timestamp 1669390400
transform -1 0 14000 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _714_
timestamp 1669390400
transform -1 0 13104 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _715_
timestamp 1669390400
transform -1 0 13104 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _716_
timestamp 1669390400
transform 1 0 9632 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _717_
timestamp 1669390400
transform 1 0 13776 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _718_
timestamp 1669390400
transform 1 0 14112 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _719_
timestamp 1669390400
transform -1 0 20944 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _720_
timestamp 1669390400
transform 1 0 17584 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _721_
timestamp 1669390400
transform 1 0 16352 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _722_
timestamp 1669390400
transform 1 0 15904 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _723_
timestamp 1669390400
transform 1 0 24080 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _724_
timestamp 1669390400
transform 1 0 19824 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _725_
timestamp 1669390400
transform -1 0 22736 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _726_
timestamp 1669390400
transform -1 0 23408 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _727_
timestamp 1669390400
transform -1 0 24416 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _728_
timestamp 1669390400
transform 1 0 26320 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _729_
timestamp 1669390400
transform 1 0 29792 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _730_
timestamp 1669390400
transform 1 0 32032 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _731_
timestamp 1669390400
transform -1 0 36736 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _732_
timestamp 1669390400
transform -1 0 36736 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _733_
timestamp 1669390400
transform 1 0 32480 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _734_
timestamp 1669390400
transform 1 0 32256 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _735_
timestamp 1669390400
transform 1 0 32144 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _736_
timestamp 1669390400
transform 1 0 33488 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _737_
timestamp 1669390400
transform 1 0 32256 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _738_
timestamp 1669390400
transform 1 0 29008 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _739_
timestamp 1669390400
transform 1 0 26880 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _740_
timestamp 1669390400
transform 1 0 25872 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _741_
timestamp 1669390400
transform 1 0 20384 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _742_
timestamp 1669390400
transform 1 0 20384 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _743_
timestamp 1669390400
transform 1 0 21504 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _744_
timestamp 1669390400
transform 1 0 17696 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 25088 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform 1 0 22848 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform -1 0 28448 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input1 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21952 0 1 3136
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 38752 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 39312 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform -1 0 40768 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform -1 0 41328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 40544 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform -1 0 40544 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform -1 0 26992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform -1 0 27216 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform -1 0 30912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 29904 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform 1 0 29456 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform -1 0 33264 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform -1 0 34832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform -1 0 35280 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform -1 0 38752 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform 1 0 1680 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18 gfth/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38752 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 3248 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform 1 0 14672 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 15344 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform 1 0 17584 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform 1 0 17472 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform 1 0 19264 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform 1 0 21504 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform -1 0 3360 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform -1 0 5152 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 5264 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 5712 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 7616 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform 1 0 7504 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform 1 0 9632 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform 1 0 11424 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform 1 0 13440 0 1 3136
box -86 -86 1654 870
<< labels >>
flabel metal3 s 43200 21952 44000 22064 0 FreeSans 448 0 0 0 bs
port 0 nsew signal tristate
flabel metal2 s 21952 43200 22064 44000 0 FreeSans 448 90 0 0 clk
port 1 nsew signal input
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 co[0]
port 2 nsew signal input
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 co[10]
port 3 nsew signal input
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 co[11]
port 4 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 co[12]
port 5 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 co[13]
port 6 nsew signal input
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 co[14]
port 7 nsew signal input
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 co[15]
port 8 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 co[1]
port 9 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 co[2]
port 10 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 co[3]
port 11 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 co[4]
port 12 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 co[5]
port 13 nsew signal input
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 co[6]
port 14 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 co[7]
port 15 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 co[8]
port 16 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 co[9]
port 17 nsew signal input
flabel metal3 s 0 21952 800 22064 0 FreeSans 448 0 0 0 st
port 18 nsew signal input
flabel metal4 s 4448 3076 4768 40828 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 35168 3076 35488 40828 0 FreeSans 1280 90 0 0 vdd
port 19 nsew power bidirectional
flabel metal4 s 19808 3076 20128 40828 0 FreeSans 1280 90 0 0 vss
port 20 nsew ground bidirectional
flabel metal2 s 1120 0 1232 800 0 FreeSans 448 90 0 0 x[0]
port 21 nsew signal tristate
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 x[10]
port 22 nsew signal tristate
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 x[11]
port 23 nsew signal tristate
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 x[12]
port 24 nsew signal tristate
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 x[13]
port 25 nsew signal tristate
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 x[14]
port 26 nsew signal tristate
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 x[15]
port 27 nsew signal tristate
flabel metal2 s 2464 0 2576 800 0 FreeSans 448 90 0 0 x[1]
port 28 nsew signal tristate
flabel metal2 s 3808 0 3920 800 0 FreeSans 448 90 0 0 x[2]
port 29 nsew signal tristate
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 x[3]
port 30 nsew signal tristate
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 x[4]
port 31 nsew signal tristate
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 x[5]
port 32 nsew signal tristate
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 x[6]
port 33 nsew signal tristate
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 x[7]
port 34 nsew signal tristate
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 x[8]
port 35 nsew signal tristate
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 x[9]
port 36 nsew signal tristate
rlabel metal1 21952 39984 21952 39984 0 vdd
rlabel metal1 21952 40768 21952 40768 0 vss
rlabel metal2 5768 12040 5768 12040 0 Datapath.i\[0\]
rlabel metal2 15400 7168 15400 7168 0 Datapath.i\[10\]
rlabel metal2 16744 15624 16744 15624 0 Datapath.i\[11\]
rlabel metal2 17864 3920 17864 3920 0 Datapath.i\[12\]
rlabel metal2 18648 8008 18648 8008 0 Datapath.i\[13\]
rlabel metal2 19432 11760 19432 11760 0 Datapath.i\[14\]
rlabel metal3 17808 9128 17808 9128 0 Datapath.i\[15\]
rlabel metal3 4480 6552 4480 6552 0 Datapath.i\[1\]
rlabel metal3 5992 6664 5992 6664 0 Datapath.i\[2\]
rlabel metal3 7616 10584 7616 10584 0 Datapath.i\[3\]
rlabel metal2 4816 12040 4816 12040 0 Datapath.i\[4\]
rlabel metal2 2856 10920 2856 10920 0 Datapath.i\[5\]
rlabel metal2 10920 11424 10920 11424 0 Datapath.i\[6\]
rlabel metal2 2296 7784 2296 7784 0 Datapath.i\[7\]
rlabel metal2 10080 10696 10080 10696 0 Datapath.i\[8\]
rlabel metal2 12936 8848 12936 8848 0 Datapath.i\[9\]
rlabel metal3 24696 10696 24696 10696 0 Datapath.k\[0\]
rlabel metal2 41832 8008 41832 8008 0 Datapath.k\[10\]
rlabel metal2 40600 11200 40600 11200 0 Datapath.k\[11\]
rlabel metal2 36344 20888 36344 20888 0 Datapath.k\[12\]
rlabel metal2 35336 16128 35336 16128 0 Datapath.k\[13\]
rlabel metal2 35448 17752 35448 17752 0 Datapath.k\[14\]
rlabel metal2 31528 17976 31528 17976 0 Datapath.k\[15\]
rlabel metal3 29736 14280 29736 14280 0 Datapath.k\[16\]
rlabel metal2 31640 17528 31640 17528 0 Datapath.k\[17\]
rlabel metal2 25480 16408 25480 16408 0 Datapath.k\[18\]
rlabel metal2 23464 17080 23464 17080 0 Datapath.k\[19\]
rlabel metal2 27608 22120 27608 22120 0 Datapath.k\[1\]
rlabel metal2 27496 21448 27496 21448 0 Datapath.k\[2\]
rlabel metal3 21504 17752 21504 17752 0 Datapath.k\[3\]
rlabel metal3 23632 20776 23632 20776 0 Datapath.k\[4\]
rlabel metal2 26824 5656 26824 5656 0 Datapath.k\[5\]
rlabel metal2 38920 21952 38920 21952 0 Datapath.k\[6\]
rlabel metal2 31864 23856 31864 23856 0 Datapath.k\[7\]
rlabel metal3 34216 17192 34216 17192 0 Datapath.k\[8\]
rlabel metal2 26264 22512 26264 22512 0 Datapath.k\[9\]
rlabel metal2 24584 14672 24584 14672 0 FSM.CS\[0\]
rlabel metal2 20776 13272 20776 13272 0 FSM.CS\[1\]
rlabel metal2 22120 14000 22120 14000 0 FSM.NS\[0\]
rlabel metal2 22792 13552 22792 13552 0 FSM.NS\[1\]
rlabel metal3 15456 8344 15456 8344 0 _000_
rlabel metal3 7840 5208 7840 5208 0 _001_
rlabel metal2 8680 7000 8680 7000 0 _002_
rlabel metal3 8400 9240 8400 9240 0 _003_
rlabel metal2 6888 11760 6888 11760 0 _004_
rlabel metal3 9632 12264 9632 12264 0 _005_
rlabel metal2 13048 10752 13048 10752 0 _006_
rlabel metal3 11816 8344 11816 8344 0 _007_
rlabel metal3 11872 6104 11872 6104 0 _008_
rlabel metal2 10584 4480 10584 4480 0 _009_
rlabel metal2 14728 6328 14728 6328 0 _010_
rlabel metal2 15736 5488 15736 5488 0 _011_
rlabel metal2 19992 4480 19992 4480 0 _012_
rlabel metal2 17024 4200 17024 4200 0 _013_
rlabel metal2 16968 10976 16968 10976 0 _014_
rlabel metal2 17024 8344 17024 8344 0 _015_
rlabel metal2 24696 10416 24696 10416 0 _016_
rlabel metal3 21672 9912 21672 9912 0 _017_
rlabel metal2 21952 8344 21952 8344 0 _018_
rlabel metal2 22456 6216 22456 6216 0 _019_
rlabel metal2 23464 5432 23464 5432 0 _020_
rlabel metal2 27720 3920 27720 3920 0 _021_
rlabel metal3 30408 4424 30408 4424 0 _022_
rlabel metal3 32144 6552 32144 6552 0 _023_
rlabel metal3 36624 5768 36624 5768 0 _024_
rlabel metal2 35896 4424 35896 4424 0 _025_
rlabel metal3 34944 8344 34944 8344 0 _026_
rlabel metal2 33208 10248 33208 10248 0 _027_
rlabel metal2 33096 13216 33096 13216 0 _028_
rlabel metal3 33600 16856 33600 16856 0 _029_
rlabel metal2 33208 16856 33208 16856 0 _030_
rlabel metal2 29848 13048 29848 13048 0 _031_
rlabel metal2 27384 16296 27384 16296 0 _032_
rlabel metal2 25984 15512 25984 15512 0 _033_
rlabel metal3 21672 15400 21672 15400 0 _034_
rlabel metal2 21784 18032 21784 18032 0 _035_
rlabel metal2 31416 22568 31416 22568 0 _036_
rlabel metal2 3192 9464 3192 9464 0 _037_
rlabel metal2 36176 20776 36176 20776 0 _038_
rlabel metal1 37688 21336 37688 21336 0 _039_
rlabel metal2 15008 15848 15008 15848 0 _040_
rlabel metal3 33768 11144 33768 11144 0 _041_
rlabel metal2 28000 21224 28000 21224 0 _042_
rlabel metal2 3192 5264 3192 5264 0 _043_
rlabel metal3 6160 6440 6160 6440 0 _044_
rlabel metal2 7448 9520 7448 9520 0 _045_
rlabel metal2 32984 24080 32984 24080 0 _046_
rlabel metal2 3192 7504 3192 7504 0 _047_
rlabel metal2 3640 4760 3640 4760 0 _048_
rlabel metal3 6160 4984 6160 4984 0 _049_
rlabel metal2 8568 10528 8568 10528 0 _050_
rlabel metal2 1960 9352 1960 9352 0 _051_
rlabel metal2 10696 8512 10696 8512 0 _052_
rlabel metal2 1848 8568 1848 8568 0 _053_
rlabel metal2 14336 4536 14336 4536 0 _054_
rlabel metal2 2240 6104 2240 6104 0 _055_
rlabel metal2 20384 17416 20384 17416 0 _056_
rlabel metal2 17752 9856 17752 9856 0 _057_
rlabel metal2 18200 11312 18200 11312 0 _058_
rlabel metal3 18480 9912 18480 9912 0 _059_
rlabel metal3 28000 21000 28000 21000 0 _060_
rlabel metal3 22400 18984 22400 18984 0 _061_
rlabel metal2 2632 6496 2632 6496 0 _062_
rlabel metal2 21672 13944 21672 13944 0 _063_
rlabel metal2 29288 20804 29288 20804 0 _064_
rlabel metal3 16968 12264 16968 12264 0 _065_
rlabel metal3 22512 13048 22512 13048 0 _066_
rlabel metal2 41776 16968 41776 16968 0 _067_
rlabel metal2 40488 17808 40488 17808 0 _068_
rlabel metal2 25256 23184 25256 23184 0 _069_
rlabel metal2 24696 3108 24696 3108 0 _070_
rlabel metal2 23800 5096 23800 5096 0 _071_
rlabel metal2 24080 6888 24080 6888 0 _072_
rlabel metal3 20440 10024 20440 10024 0 _073_
rlabel metal2 22568 12712 22568 12712 0 _074_
rlabel metal3 40992 23240 40992 23240 0 _075_
rlabel metal2 37576 6160 37576 6160 0 _076_
rlabel metal2 42056 15680 42056 15680 0 _077_
rlabel metal3 31080 12152 31080 12152 0 _078_
rlabel metal2 40488 9856 40488 9856 0 _079_
rlabel metal3 41160 9128 41160 9128 0 _080_
rlabel metal2 41048 22008 41048 22008 0 _081_
rlabel metal2 30576 15848 30576 15848 0 _082_
rlabel metal3 29904 18200 29904 18200 0 _083_
rlabel metal3 29960 15848 29960 15848 0 _084_
rlabel metal2 30632 12600 30632 12600 0 _085_
rlabel metal2 25928 12488 25928 12488 0 _086_
rlabel metal3 27776 9800 27776 9800 0 _087_
rlabel metal2 33880 15512 33880 15512 0 _088_
rlabel metal3 32704 16072 32704 16072 0 _089_
rlabel metal2 27496 19600 27496 19600 0 _090_
rlabel metal3 27160 12824 27160 12824 0 _091_
rlabel metal2 26432 9576 26432 9576 0 _092_
rlabel metal2 36792 20804 36792 20804 0 _093_
rlabel metal2 37240 18088 37240 18088 0 _094_
rlabel metal2 23016 6384 23016 6384 0 _095_
rlabel metal3 28056 21336 28056 21336 0 _096_
rlabel metal3 37464 15288 37464 15288 0 _097_
rlabel metal2 34888 15232 34888 15232 0 _098_
rlabel metal2 37576 13384 37576 13384 0 _099_
rlabel metal2 28392 20440 28392 20440 0 _100_
rlabel metal2 26600 9800 26600 9800 0 _101_
rlabel metal3 2632 6104 2632 6104 0 _102_
rlabel metal2 35896 22512 35896 22512 0 _103_
rlabel metal2 26712 9576 26712 9576 0 _104_
rlabel metal2 14616 10192 14616 10192 0 _105_
rlabel metal3 6888 8008 6888 8008 0 _106_
rlabel metal2 6328 6440 6328 6440 0 _107_
rlabel metal3 5880 6104 5880 6104 0 _108_
rlabel metal3 5376 7560 5376 7560 0 _109_
rlabel metal2 6160 9128 6160 9128 0 _110_
rlabel metal2 4928 8008 4928 8008 0 _111_
rlabel metal2 6776 7728 6776 7728 0 _112_
rlabel metal3 7056 9016 7056 9016 0 _113_
rlabel metal2 8232 9688 8232 9688 0 _114_
rlabel metal2 7560 9800 7560 9800 0 _115_
rlabel metal2 7448 11368 7448 11368 0 _116_
rlabel metal3 7392 11256 7392 11256 0 _117_
rlabel metal2 6776 11200 6776 11200 0 _118_
rlabel metal2 9912 11704 9912 11704 0 _119_
rlabel metal3 26712 22232 26712 22232 0 _120_
rlabel metal2 2744 6160 2744 6160 0 _121_
rlabel metal3 8008 9128 8008 9128 0 _122_
rlabel metal2 10584 9688 10584 9688 0 _123_
rlabel metal2 10528 12152 10528 12152 0 _124_
rlabel metal3 10696 11144 10696 11144 0 _125_
rlabel metal2 11872 11480 11872 11480 0 _126_
rlabel metal2 11144 11592 11144 11592 0 _127_
rlabel metal2 2408 7532 2408 7532 0 _128_
rlabel metal2 12824 12432 12824 12432 0 _129_
rlabel metal2 11816 10304 11816 10304 0 _130_
rlabel metal2 6440 13440 6440 13440 0 _131_
rlabel metal2 11144 6608 11144 6608 0 _132_
rlabel metal3 11704 4984 11704 4984 0 _133_
rlabel metal2 14840 7112 14840 7112 0 _134_
rlabel metal2 8904 7616 8904 7616 0 _135_
rlabel metal2 4312 8120 4312 8120 0 _136_
rlabel metal3 7560 7448 7560 7448 0 _137_
rlabel metal2 1848 5208 1848 5208 0 _138_
rlabel metal2 14840 11984 14840 11984 0 _139_
rlabel metal2 15512 8176 15512 8176 0 _140_
rlabel metal2 16296 16240 16296 16240 0 _141_
rlabel metal2 17416 7616 17416 7616 0 _142_
rlabel metal2 2520 7616 2520 7616 0 _143_
rlabel metal2 13608 8960 13608 8960 0 _144_
rlabel metal2 19376 6664 19376 6664 0 _145_
rlabel metal2 17584 15848 17584 15848 0 _146_
rlabel metal3 18424 16856 18424 16856 0 _147_
rlabel metal2 19936 5096 19936 5096 0 _148_
rlabel metal2 18984 6160 18984 6160 0 _149_
rlabel metal2 16856 4984 16856 4984 0 _150_
rlabel metal2 16856 10864 16856 10864 0 _151_
rlabel metal2 18256 9240 18256 9240 0 _152_
rlabel metal3 17752 8904 17752 8904 0 _153_
rlabel metal3 18312 9800 18312 9800 0 _154_
rlabel metal3 26656 13720 26656 13720 0 _155_
rlabel metal3 25200 13608 25200 13608 0 _156_
rlabel metal2 24808 12040 24808 12040 0 _157_
rlabel metal2 30520 24360 30520 24360 0 _158_
rlabel metal2 16632 6552 16632 6552 0 _159_
rlabel metal2 23128 7840 23128 7840 0 _160_
rlabel metal3 29904 10696 29904 10696 0 _161_
rlabel metal3 26824 19992 26824 19992 0 _162_
rlabel metal2 25816 11816 25816 11816 0 _163_
rlabel metal2 25032 9912 25032 9912 0 _164_
rlabel metal3 26544 21560 26544 21560 0 _165_
rlabel metal2 22344 8680 22344 8680 0 _166_
rlabel metal2 27160 9296 27160 9296 0 _167_
rlabel metal3 26488 20776 26488 20776 0 _168_
rlabel metal2 23576 9408 23576 9408 0 _169_
rlabel metal3 26376 20104 26376 20104 0 _170_
rlabel metal3 24808 9688 24808 9688 0 _171_
rlabel metal2 23296 6664 23296 6664 0 _172_
rlabel metal2 23688 6384 23688 6384 0 _173_
rlabel metal3 23856 9016 23856 9016 0 _174_
rlabel metal2 27944 20496 27944 20496 0 _175_
rlabel metal3 14616 3304 14616 3304 0 _176_
rlabel metal2 25032 6048 25032 6048 0 _177_
rlabel metal2 29400 22456 29400 22456 0 _178_
rlabel metal3 27496 18704 27496 18704 0 _179_
rlabel metal2 26824 8120 26824 8120 0 _180_
rlabel metal2 28840 22120 28840 22120 0 _181_
rlabel metal2 25704 7784 25704 7784 0 _182_
rlabel metal2 25984 6104 25984 6104 0 _183_
rlabel metal3 30520 6664 30520 6664 0 _184_
rlabel metal2 28616 22960 28616 22960 0 _185_
rlabel metal2 26936 22008 26936 22008 0 _186_
rlabel metal3 32256 7448 32256 7448 0 _187_
rlabel metal2 31752 22848 31752 22848 0 _188_
rlabel metal2 27720 6944 27720 6944 0 _189_
rlabel metal2 27832 4144 27832 4144 0 _190_
rlabel metal2 28056 3864 28056 3864 0 _191_
rlabel metal2 26712 6160 26712 6160 0 _192_
rlabel metal2 27664 6104 27664 6104 0 _193_
rlabel metal2 30128 22456 30128 22456 0 _194_
rlabel metal2 41384 20440 41384 20440 0 _195_
rlabel metal2 32200 10360 32200 10360 0 _196_
rlabel metal2 31752 8456 31752 8456 0 _197_
rlabel metal2 30968 22008 30968 22008 0 _198_
rlabel metal2 31192 9800 31192 9800 0 _199_
rlabel metal2 32200 22848 32200 22848 0 _200_
rlabel metal2 30184 8120 30184 8120 0 _201_
rlabel metal2 30912 6104 30912 6104 0 _202_
rlabel metal2 38416 17192 38416 17192 0 _203_
rlabel metal3 34832 20216 34832 20216 0 _204_
rlabel metal2 36680 17136 36680 17136 0 _205_
rlabel metal3 35504 18200 35504 18200 0 _206_
rlabel metal2 32648 21112 32648 21112 0 _207_
rlabel metal2 31808 9240 31808 9240 0 _208_
rlabel metal2 33096 24528 33096 24528 0 _209_
rlabel metal3 31864 9016 31864 9016 0 _210_
rlabel metal2 31472 6664 31472 6664 0 _211_
rlabel metal2 31696 6664 31696 6664 0 _212_
rlabel metal3 36904 23520 36904 23520 0 _213_
rlabel metal3 31528 22344 31528 22344 0 _214_
rlabel metal3 29400 22568 29400 22568 0 _215_
rlabel metal2 29736 10080 29736 10080 0 _216_
rlabel metal3 39648 23016 39648 23016 0 _217_
rlabel metal2 28728 7168 28728 7168 0 _218_
rlabel metal2 31080 20804 31080 20804 0 _219_
rlabel metal2 40432 21448 40432 21448 0 _220_
rlabel metal3 41272 8120 41272 8120 0 _221_
rlabel metal3 40656 10808 40656 10808 0 _222_
rlabel metal3 41384 12376 41384 12376 0 _223_
rlabel metal4 41720 14896 41720 14896 0 _224_
rlabel metal2 41832 11312 41832 11312 0 _225_
rlabel metal2 41944 17808 41944 17808 0 _226_
rlabel metal2 42112 21784 42112 21784 0 _227_
rlabel metal4 39368 8512 39368 8512 0 _228_
rlabel metal2 37352 6272 37352 6272 0 _229_
rlabel metal3 34888 3304 34888 3304 0 _230_
rlabel metal2 24136 21392 24136 21392 0 _231_
rlabel metal2 41496 13720 41496 13720 0 _232_
rlabel metal3 41384 19320 41384 19320 0 _233_
rlabel metal2 24808 23128 24808 23128 0 _234_
rlabel metal3 40264 3528 40264 3528 0 _235_
rlabel metal3 41496 3192 41496 3192 0 _236_
rlabel metal2 36680 7168 36680 7168 0 _237_
rlabel metal2 39256 7112 39256 7112 0 _238_
rlabel metal2 41888 7560 41888 7560 0 _239_
rlabel metal2 39816 6496 39816 6496 0 _240_
rlabel metal2 41104 6552 41104 6552 0 _241_
rlabel metal3 41160 9576 41160 9576 0 _242_
rlabel metal2 41272 5768 41272 5768 0 _243_
rlabel metal2 38024 9744 38024 9744 0 _244_
rlabel metal2 38584 6384 38584 6384 0 _245_
rlabel metal3 37128 8008 37128 8008 0 _246_
rlabel metal2 35840 7672 35840 7672 0 _247_
rlabel metal2 40936 9968 40936 9968 0 _248_
rlabel metal2 38696 10192 38696 10192 0 _249_
rlabel metal2 40488 12208 40488 12208 0 _250_
rlabel metal2 40376 11424 40376 11424 0 _251_
rlabel metal3 37464 10528 37464 10528 0 _252_
rlabel metal3 34832 10472 34832 10472 0 _253_
rlabel metal3 33488 10808 33488 10808 0 _254_
rlabel metal2 40824 10304 40824 10304 0 _255_
rlabel metal2 41608 7336 41608 7336 0 _256_
rlabel metal2 39704 12544 39704 12544 0 _257_
rlabel metal3 41552 7224 41552 7224 0 _258_
rlabel metal2 39256 11284 39256 11284 0 _259_
rlabel metal3 41384 12712 41384 12712 0 _260_
rlabel metal2 38808 12376 38808 12376 0 _261_
rlabel metal3 39480 12824 39480 12824 0 _262_
rlabel metal3 40264 11592 40264 11592 0 _263_
rlabel metal2 38472 12936 38472 12936 0 _264_
rlabel metal2 39704 13384 39704 13384 0 _265_
rlabel metal3 39816 12264 39816 12264 0 _266_
rlabel metal2 34160 13720 34160 13720 0 _267_
rlabel metal2 35560 13048 35560 13048 0 _268_
rlabel metal2 40488 15736 40488 15736 0 _269_
rlabel metal3 36624 13832 36624 13832 0 _270_
rlabel metal3 36456 12824 36456 12824 0 _271_
rlabel metal3 37576 13496 37576 13496 0 _272_
rlabel metal2 36624 13944 36624 13944 0 _273_
rlabel metal2 36288 13944 36288 13944 0 _274_
rlabel metal3 34440 14504 34440 14504 0 _275_
rlabel metal2 32928 14504 32928 14504 0 _276_
rlabel metal2 38920 14000 38920 14000 0 _277_
rlabel metal2 38584 15624 38584 15624 0 _278_
rlabel metal2 38920 15064 38920 15064 0 _279_
rlabel metal2 39032 17136 39032 17136 0 _280_
rlabel metal2 39760 15512 39760 15512 0 _281_
rlabel metal2 35896 15680 35896 15680 0 _282_
rlabel metal2 36008 17584 36008 17584 0 _283_
rlabel metal3 37352 16968 37352 16968 0 _284_
rlabel metal3 40096 16856 40096 16856 0 _285_
rlabel metal2 38248 17304 38248 17304 0 _286_
rlabel metal2 38808 16912 38808 16912 0 _287_
rlabel metal2 33096 16744 33096 16744 0 _288_
rlabel metal3 33544 16184 33544 16184 0 _289_
rlabel metal3 38024 17080 38024 17080 0 _290_
rlabel metal3 36848 17080 36848 17080 0 _291_
rlabel metal2 36344 15624 36344 15624 0 _292_
rlabel metal2 37464 15848 37464 15848 0 _293_
rlabel metal2 37688 17136 37688 17136 0 _294_
rlabel metal3 36904 15960 36904 15960 0 _295_
rlabel metal3 37016 16072 37016 16072 0 _296_
rlabel metal3 37352 15848 37352 15848 0 _297_
rlabel metal2 29512 12656 29512 12656 0 _298_
rlabel metal3 29456 12936 29456 12936 0 _299_
rlabel metal2 38696 15848 38696 15848 0 _300_
rlabel metal3 39368 14392 39368 14392 0 _301_
rlabel metal2 40768 14392 40768 14392 0 _302_
rlabel metal4 39816 11200 39816 11200 0 _303_
rlabel metal2 31528 15736 31528 15736 0 _304_
rlabel metal2 40376 14952 40376 14952 0 _305_
rlabel metal3 37912 15400 37912 15400 0 _306_
rlabel metal3 39536 15288 39536 15288 0 _307_
rlabel metal2 31304 16352 31304 16352 0 _308_
rlabel metal2 31640 15848 31640 15848 0 _309_
rlabel metal3 33040 15288 33040 15288 0 _310_
rlabel metal3 30520 15288 30520 15288 0 _311_
rlabel metal3 33208 15176 33208 15176 0 _312_
rlabel metal3 30016 14728 30016 14728 0 _313_
rlabel metal3 31416 16072 31416 16072 0 _314_
rlabel metal3 31024 15512 31024 15512 0 _315_
rlabel metal4 27384 16688 27384 16688 0 _316_
rlabel metal3 24472 19208 24472 19208 0 _317_
rlabel metal2 27272 15624 27272 15624 0 _318_
rlabel metal2 27496 16296 27496 16296 0 _319_
rlabel metal3 30016 15512 30016 15512 0 _320_
rlabel metal2 30408 17584 30408 17584 0 _321_
rlabel metal2 26936 15568 26936 15568 0 _322_
rlabel metal2 29960 15960 29960 15960 0 _323_
rlabel metal3 28448 15288 28448 15288 0 _324_
rlabel metal3 26432 15288 26432 15288 0 _325_
rlabel metal2 25592 15568 25592 15568 0 _326_
rlabel metal2 30856 17080 30856 17080 0 _327_
rlabel metal3 30744 17416 30744 17416 0 _328_
rlabel metal3 28504 17752 28504 17752 0 _329_
rlabel metal2 26264 17248 26264 17248 0 _330_
rlabel metal2 24808 17752 24808 17752 0 _331_
rlabel metal3 27216 17528 27216 17528 0 _332_
rlabel metal3 26600 17864 26600 17864 0 _333_
rlabel metal2 25480 18424 25480 18424 0 _334_
rlabel metal3 25480 19096 25480 19096 0 _335_
rlabel metal2 22008 16632 22008 16632 0 _336_
rlabel metal2 22344 16128 22344 16128 0 _337_
rlabel metal2 23912 16184 23912 16184 0 _338_
rlabel metal2 24136 17696 24136 17696 0 _339_
rlabel metal2 23464 17976 23464 17976 0 _340_
rlabel metal2 21952 17640 21952 17640 0 _341_
rlabel metal2 21672 18144 21672 18144 0 _342_
rlabel metal2 23128 17360 23128 17360 0 _343_
rlabel metal2 40040 22120 40040 22120 0 bs
rlabel metal2 22008 41146 22008 41146 0 clk
rlabel metal2 16632 15176 16632 15176 0 clknet_0_clk
rlabel metal2 3080 7952 3080 7952 0 clknet_2_0__leaf_clk
rlabel metal2 19712 15848 19712 15848 0 clknet_2_1__leaf_clk
rlabel metal2 25592 22736 25592 22736 0 clknet_2_2__leaf_clk
rlabel metal2 29512 18704 29512 18704 0 clknet_2_3__leaf_clk
rlabel metal3 13104 2968 13104 2968 0 co[0]
rlabel metal3 42280 23016 42280 23016 0 co[10]
rlabel metal3 41216 23800 41216 23800 0 co[11]
rlabel metal3 22568 3080 22568 3080 0 co[12]
rlabel metal2 40152 1918 40152 1918 0 co[13]
rlabel metal2 41384 3080 41384 3080 0 co[14]
rlabel metal3 40320 23576 40320 23576 0 co[15]
rlabel metal2 19488 17416 19488 17416 0 co[1]
rlabel metal2 25368 1974 25368 1974 0 co[2]
rlabel metal3 24024 21448 24024 21448 0 co[3]
rlabel metal3 23240 24024 23240 24024 0 co[4]
rlabel metal2 1624 11760 1624 11760 0 co[5]
rlabel metal3 32984 23688 32984 23688 0 co[6]
rlabel metal3 41664 22120 41664 22120 0 co[7]
rlabel metal3 38528 23912 38528 23912 0 co[8]
rlabel metal2 1736 10360 1736 10360 0 co[9]
rlabel metal2 25256 20356 25256 20356 0 net1
rlabel metal2 24192 5096 24192 5096 0 net10
rlabel metal2 26152 5600 26152 5600 0 net11
rlabel metal3 31640 5208 31640 5208 0 net12
rlabel metal3 31976 5880 31976 5880 0 net13
rlabel metal3 32928 5656 32928 5656 0 net14
rlabel metal2 32760 4592 32760 4592 0 net15
rlabel metal3 36680 5096 36680 5096 0 net16
rlabel metal2 3360 22456 3360 22456 0 net17
rlabel metal2 38416 22232 38416 22232 0 net18
rlabel metal2 2968 4760 2968 4760 0 net19
rlabel metal3 35336 5096 35336 5096 0 net2
rlabel metal2 14840 10696 14840 10696 0 net20
rlabel metal3 15400 16856 15400 16856 0 net21
rlabel metal2 2184 5432 2184 5432 0 net22
rlabel metal2 14168 5768 14168 5768 0 net23
rlabel metal2 17976 9576 17976 9576 0 net24
rlabel metal2 21784 6496 21784 6496 0 net25
rlabel metal2 3080 4200 3080 4200 0 net26
rlabel metal2 4536 3528 4536 3528 0 net27
rlabel metal2 4872 5880 4872 5880 0 net28
rlabel metal3 4928 4424 4928 4424 0 net29
rlabel metal4 35896 7336 35896 7336 0 net3
rlabel metal3 6384 4872 6384 4872 0 net30
rlabel metal2 7896 4592 7896 4592 0 net31
rlabel metal3 7336 3528 7336 3528 0 net32
rlabel metal2 11312 3528 11312 3528 0 net33
rlabel metal2 13608 3976 13608 3976 0 net34
rlabel metal2 36848 21672 36848 21672 0 net4
rlabel metal2 23464 21000 23464 21000 0 net5
rlabel metal2 22568 19712 22568 19712 0 net6
rlabel metal3 31080 20552 31080 20552 0 net7
rlabel metal3 24024 16968 24024 16968 0 net8
rlabel metal2 23968 5096 23968 5096 0 net9
rlabel metal2 1848 21896 1848 21896 0 st
rlabel metal2 1176 2478 1176 2478 0 x[0]
rlabel metal2 14616 2478 14616 2478 0 x[10]
rlabel metal2 15960 2058 15960 2058 0 x[11]
rlabel metal3 17864 5208 17864 5208 0 x[12]
rlabel metal2 18648 2198 18648 2198 0 x[13]
rlabel metal2 19992 1862 19992 1862 0 x[14]
rlabel metal3 21840 3976 21840 3976 0 x[15]
rlabel metal2 2520 2198 2520 2198 0 x[1]
rlabel metal2 3864 2086 3864 2086 0 x[2]
rlabel metal3 5656 4200 5656 4200 0 x[3]
rlabel metal2 6552 2198 6552 2198 0 x[4]
rlabel metal2 7896 854 7896 854 0 x[5]
rlabel metal2 9240 2058 9240 2058 0 x[6]
rlabel metal2 10584 2198 10584 2198 0 x[7]
rlabel metal2 11928 2058 11928 2058 0 x[8]
rlabel metal3 13776 3640 13776 3640 0 x[9]
<< properties >>
string FIXED_BBOX 0 0 44000 44000
<< end >>
